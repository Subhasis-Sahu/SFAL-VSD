# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o311ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.775000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.055000 3.615000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 1.055000 5.885000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 1.055000 7.695000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.865000 1.055000 9.090000 1.315000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.241000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055000 1.485000 9.575000 1.725000 ;
        RECT 4.055000 1.725000 4.305000 2.115000 ;
        RECT 4.975000 1.725000 5.145000 2.115000 ;
        RECT 5.815000 1.725000 6.005000 2.465000 ;
        RECT 6.675000 1.725000 6.845000 2.465000 ;
        RECT 7.515000 1.725000 7.685000 2.465000 ;
        RECT 7.895000 0.655000 9.575000 0.885000 ;
        RECT 8.355000 1.725000 8.525000 2.465000 ;
        RECT 9.195000 1.725000 9.575000 2.465000 ;
        RECT 9.260000 0.885000 9.575000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.085000  0.085000 0.505000 0.885000 ;
        RECT 1.015000  0.085000 1.345000 0.485000 ;
        RECT 1.855000  0.085000 2.185000 0.485000 ;
        RECT 2.695000  0.085000 3.025000 0.485000 ;
        RECT 3.535000  0.085000 3.885000 0.485000 ;
        RECT 4.395000  0.085000 4.725000 0.485000 ;
        RECT 5.235000  0.085000 5.585000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.595000 1.895000 0.925000 2.635000 ;
        RECT 1.435000 1.895000 1.765000 2.635000 ;
        RECT 6.175000 1.895000 6.505000 2.635000 ;
        RECT 7.015000 1.895000 7.345000 2.635000 ;
        RECT 7.855000 1.895000 8.185000 2.635000 ;
        RECT 8.695000 1.895000 9.025000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.485000 3.865000 1.725000 ;
      RECT 0.085000 1.725000 0.405000 2.465000 ;
      RECT 0.675000 0.255000 0.845000 0.655000 ;
      RECT 0.675000 0.655000 7.385000 0.885000 ;
      RECT 1.095000 1.725000 1.265000 2.465000 ;
      RECT 1.515000 0.255000 1.685000 0.655000 ;
      RECT 1.935000 1.725000 2.105000 2.465000 ;
      RECT 2.275000 1.895000 2.605000 2.295000 ;
      RECT 2.275000 2.295000 5.645000 2.465000 ;
      RECT 2.355000 0.255000 2.525000 0.655000 ;
      RECT 2.775000 1.725000 2.945000 2.115000 ;
      RECT 3.115000 1.895000 3.445000 2.295000 ;
      RECT 3.195000 0.255000 3.365000 0.655000 ;
      RECT 3.615000 1.725000 3.865000 2.115000 ;
      RECT 4.055000 0.255000 4.225000 0.655000 ;
      RECT 4.475000 1.895000 4.805000 2.295000 ;
      RECT 4.895000 0.255000 5.065000 0.655000 ;
      RECT 5.315000 1.895000 5.645000 2.295000 ;
      RECT 5.755000 0.255000 9.575000 0.485000 ;
      RECT 7.555000 0.485000 7.725000 0.885000 ;
  END
END sky130_fd_sc_hd__o311ai_4
END LIBRARY
