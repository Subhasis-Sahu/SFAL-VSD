# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__or4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235000 0.995000 3.405000 1.445000 ;
        RECT 3.235000 1.445000 3.670000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 0.995000 3.005000 1.450000 ;
        RECT 2.795000 1.450000 3.005000 1.785000 ;
        RECT 2.795000 1.785000 3.115000 2.375000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 1.455000 5.435000 1.625000 ;
        RECT 3.875000 1.625000 4.125000 2.465000 ;
        RECT 3.915000 0.255000 4.165000 0.725000 ;
        RECT 3.915000 0.725000 5.435000 0.905000 ;
        RECT 4.675000 0.255000 5.005000 0.725000 ;
        RECT 4.715000 1.625000 4.965000 2.465000 ;
        RECT 5.205000 0.905000 5.435000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.655000  0.085000 0.825000 0.825000 ;
        RECT 1.515000  0.085000 1.845000 0.480000 ;
        RECT 2.465000  0.085000 2.795000 0.485000 ;
        RECT 3.355000  0.085000 3.735000 0.485000 ;
        RECT 4.335000  0.085000 4.505000 0.555000 ;
        RECT 5.175000  0.085000 5.345000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.515000 2.205000 0.845000 2.635000 ;
        RECT 3.400000 1.795000 3.650000 2.635000 ;
        RECT 4.295000 1.795000 4.545000 2.635000 ;
        RECT 5.135000 1.795000 5.385000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.450000 0.400000 0.825000 ;
      RECT 0.085000 0.825000 0.255000 1.865000 ;
      RECT 0.085000 1.865000 1.295000 2.035000 ;
      RECT 0.085000 2.035000 0.345000 2.455000 ;
      RECT 0.990000 1.525000 1.595000 1.695000 ;
      RECT 1.075000 0.450000 1.245000 0.655000 ;
      RECT 1.075000 0.655000 1.595000 0.825000 ;
      RECT 1.125000 2.035000 1.295000 2.295000 ;
      RECT 1.125000 2.295000 2.445000 2.465000 ;
      RECT 1.405000 0.825000 1.595000 0.995000 ;
      RECT 1.405000 0.995000 1.695000 1.325000 ;
      RECT 1.405000 1.325000 1.595000 1.525000 ;
      RECT 1.510000 1.955000 2.105000 2.125000 ;
      RECT 1.935000 0.655000 3.745000 0.825000 ;
      RECT 1.935000 0.825000 2.105000 1.955000 ;
      RECT 2.095000 0.305000 2.265000 0.655000 ;
      RECT 2.275000 0.995000 2.445000 2.295000 ;
      RECT 2.965000 0.305000 3.135000 0.655000 ;
      RECT 3.575000 0.825000 3.745000 1.075000 ;
      RECT 3.575000 1.075000 5.035000 1.245000 ;
  END
END sky130_fd_sc_hd__or4bb_4
END LIBRARY
