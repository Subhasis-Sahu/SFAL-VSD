# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__fah_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.440000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 2.495000 1.275000 ;
        RECT 1.990000 1.275000 2.190000 1.410000 ;
        RECT 2.015000 1.410000 2.190000 1.725000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.675000 0.995000 5.925000 1.325000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.930000 1.075000 2.220000 1.120000 ;
        RECT 1.930000 1.120000 5.910000 1.260000 ;
        RECT 1.930000 1.260000 2.220000 1.305000 ;
        RECT 5.620000 1.075000 5.910000 1.120000 ;
        RECT 5.620000 1.260000 5.910000 1.305000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.475000 1.075000  9.865000 1.325000 ;
        RECT 9.690000 0.735000 10.010000 0.935000 ;
        RECT 9.690000 0.935000  9.865000 1.075000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.870000 0.270000 11.310000 0.825000 ;
        RECT 10.870000 0.825000 11.040000 1.495000 ;
        RECT 10.870000 1.495000 11.390000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.506000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.980000 0.255000 12.335000 0.825000 ;
        RECT 11.985000 1.785000 12.335000 2.465000 ;
        RECT 12.110000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.420000 0.085000 ;
        RECT  0.595000  0.085000  0.765000 0.545000 ;
        RECT  2.010000  0.085000  2.180000 0.545000 ;
        RECT  9.905000  0.085000 10.075000 0.565000 ;
        RECT 11.480000  0.085000 11.810000 0.825000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 12.420000 2.805000 ;
        RECT  0.565000 2.260000  0.930000 2.635000 ;
        RECT  2.065000 2.235000  2.395000 2.635000 ;
        RECT  9.840000 2.275000 10.175000 2.635000 ;
        RECT 11.560000 1.785000 11.815000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.255000  0.425000 0.805000 ;
      RECT  0.085000 0.805000  0.255000 1.500000 ;
      RECT  0.085000 1.500000  0.445000 1.895000 ;
      RECT  0.085000 1.895000  2.805000 2.065000 ;
      RECT  0.085000 2.065000  0.395000 2.465000 ;
      RECT  0.425000 0.995000  0.780000 1.325000 ;
      RECT  0.595000 0.735000  1.320000 0.905000 ;
      RECT  0.595000 0.905000  0.780000 0.995000 ;
      RECT  0.610000 1.325000  0.780000 1.380000 ;
      RECT  0.610000 1.380000  0.815000 1.445000 ;
      RECT  0.610000 1.445000  1.315000 1.455000 ;
      RECT  0.615000 1.455000  1.315000 1.615000 ;
      RECT  0.985000 1.615000  1.315000 1.715000 ;
      RECT  0.990000 0.255000  1.320000 0.735000 ;
      RECT  1.490000 1.445000  1.820000 1.500000 ;
      RECT  1.490000 1.500000  1.840000 1.725000 ;
      RECT  1.500000 0.255000  1.840000 0.715000 ;
      RECT  1.500000 0.715000  2.520000 0.885000 ;
      RECT  1.500000 0.885000  1.820000 0.905000 ;
      RECT  1.615000 0.905000  1.820000 1.445000 ;
      RECT  2.350000 0.255000  4.840000 0.425000 ;
      RECT  2.350000 0.425000  2.520000 0.715000 ;
      RECT  2.360000 1.445000  2.860000 1.715000 ;
      RECT  2.635000 2.065000  2.805000 2.295000 ;
      RECT  2.635000 2.295000  4.950000 2.465000 ;
      RECT  2.690000 0.595000  2.860000 1.445000 ;
      RECT  3.030000 0.425000  4.840000 0.465000 ;
      RECT  3.030000 0.465000  3.200000 1.955000 ;
      RECT  3.030000 1.955000  4.320000 2.125000 ;
      RECT  3.370000 0.635000  3.900000 0.805000 ;
      RECT  3.370000 0.805000  3.540000 1.455000 ;
      RECT  3.370000 1.455000  3.815000 1.785000 ;
      RECT  3.985000 1.785000  4.320000 1.955000 ;
      RECT  4.070000 0.645000  4.400000 0.735000 ;
      RECT  4.070000 0.735000  4.560000 0.755000 ;
      RECT  4.070000 0.755000  5.170000 0.780000 ;
      RECT  4.070000 0.780000  5.155000 0.805000 ;
      RECT  4.070000 0.805000  5.145000 0.905000 ;
      RECT  4.070000 1.075000  4.400000 1.160000 ;
      RECT  4.070000 1.160000  4.535000 1.615000 ;
      RECT  4.480000 0.905000  5.145000 0.925000 ;
      RECT  4.650000 0.465000  4.840000 0.585000 ;
      RECT  4.705000 0.925000  4.875000 2.295000 ;
      RECT  4.925000 0.735000  5.180000 0.740000 ;
      RECT  4.925000 0.740000  5.170000 0.755000 ;
      RECT  4.950000 0.715000  5.180000 0.735000 ;
      RECT  4.980000 0.690000  5.180000 0.715000 ;
      RECT  5.000000 0.655000  5.180000 0.690000 ;
      RECT  5.010000 0.255000  6.100000 0.425000 ;
      RECT  5.010000 0.425000  5.180000 0.655000 ;
      RECT  5.125000 1.150000  5.505000 1.320000 ;
      RECT  5.125000 1.320000  5.295000 2.295000 ;
      RECT  5.125000 2.295000  7.560000 2.465000 ;
      RECT  5.320000 0.865000  5.520000 0.925000 ;
      RECT  5.320000 0.925000  5.505000 1.150000 ;
      RECT  5.335000 0.840000  5.520000 0.865000 ;
      RECT  5.350000 0.595000  5.520000 0.840000 ;
      RECT  5.475000 1.700000  5.875000 2.030000 ;
      RECT  5.750000 0.425000  6.100000 0.565000 ;
      RECT  6.105000 0.740000  6.435000 1.275000 ;
      RECT  6.105000 1.445000  6.460000 1.615000 ;
      RECT  6.270000 0.255000  9.735000 0.425000 ;
      RECT  6.270000 0.425000  6.600000 0.570000 ;
      RECT  6.290000 1.615000  6.460000 1.955000 ;
      RECT  6.290000 1.955000  7.220000 2.125000 ;
      RECT  6.610000 0.755000  6.940000 0.925000 ;
      RECT  6.610000 0.925000  6.880000 1.275000 ;
      RECT  6.710000 1.275000  6.880000 1.785000 ;
      RECT  6.770000 0.595000  6.940000 0.755000 ;
      RECT  7.050000 1.060000  7.280000 1.130000 ;
      RECT  7.050000 1.130000  7.245000 1.175000 ;
      RECT  7.050000 1.175000  7.220000 1.955000 ;
      RECT  7.065000 1.045000  7.280000 1.060000 ;
      RECT  7.090000 1.010000  7.280000 1.045000 ;
      RECT  7.110000 0.595000  7.445000 0.765000 ;
      RECT  7.110000 0.765000  7.280000 1.010000 ;
      RECT  7.390000 1.275000  7.620000 1.375000 ;
      RECT  7.390000 1.375000  7.595000 1.400000 ;
      RECT  7.390000 1.400000  7.575000 1.425000 ;
      RECT  7.390000 1.425000  7.560000 2.295000 ;
      RECT  7.450000 0.995000  7.620000 1.275000 ;
      RECT  7.705000 0.425000  7.960000 0.825000 ;
      RECT  7.730000 1.510000  7.960000 2.295000 ;
      RECT  7.730000 2.295000  9.655000 2.465000 ;
      RECT  7.790000 0.825000  7.960000 1.510000 ;
      RECT  8.145000 1.955000  9.250000 2.125000 ;
      RECT  8.155000 0.595000  8.405000 0.925000 ;
      RECT  8.225000 0.925000  8.405000 1.445000 ;
      RECT  8.225000 1.445000  8.910000 1.785000 ;
      RECT  8.575000 0.595000  8.745000 1.105000 ;
      RECT  8.575000 1.105000  9.250000 1.275000 ;
      RECT  8.920000 0.685000  9.300000 0.935000 ;
      RECT  9.080000 1.275000  9.250000 1.955000 ;
      RECT  9.400000 0.425000  9.735000 0.515000 ;
      RECT  9.420000 1.495000 10.350000 1.705000 ;
      RECT  9.420000 1.705000  9.655000 2.295000 ;
      RECT 10.180000 0.995000 10.350000 1.495000 ;
      RECT 10.245000 0.285000 10.690000 0.825000 ;
      RECT 10.345000 1.875000 10.690000 2.465000 ;
      RECT 10.520000 0.825000 10.690000 1.875000 ;
      RECT 11.210000 0.995000 11.460000 1.325000 ;
      RECT 11.630000 0.995000 11.940000 1.615000 ;
    LAYER mcon ;
      RECT  2.450000 1.445000  2.620000 1.615000 ;
      RECT  3.370000 0.765000  3.540000 0.935000 ;
      RECT  3.985000 1.785000  4.155000 1.955000 ;
      RECT  4.365000 1.445000  4.535000 1.615000 ;
      RECT  5.570000 1.785000  5.740000 1.955000 ;
      RECT  6.150000 0.765000  6.320000 0.935000 ;
      RECT  6.150000 1.445000  6.320000 1.615000 ;
      RECT  6.610000 1.105000  6.780000 1.275000 ;
      RECT  8.460000 1.445000  8.630000 1.615000 ;
      RECT  8.920000 0.765000  9.090000 0.935000 ;
      RECT  9.080000 1.785000  9.250000 1.955000 ;
      RECT 10.520000 1.785000 10.690000 1.955000 ;
      RECT 11.220000 1.105000 11.390000 1.275000 ;
      RECT 11.680000 1.445000 11.850000 1.615000 ;
    LAYER met1 ;
      RECT  2.390000 1.415000  2.680000 1.460000 ;
      RECT  2.390000 1.460000  6.380000 1.600000 ;
      RECT  2.390000 1.600000  2.680000 1.645000 ;
      RECT  3.310000 0.735000  3.600000 0.780000 ;
      RECT  3.310000 0.780000  9.150000 0.920000 ;
      RECT  3.310000 0.920000  3.600000 0.965000 ;
      RECT  3.925000 1.755000  4.215000 1.800000 ;
      RECT  3.925000 1.800000  5.800000 1.940000 ;
      RECT  3.925000 1.940000  4.215000 1.985000 ;
      RECT  4.305000 1.415000  4.595000 1.460000 ;
      RECT  4.305000 1.600000  4.595000 1.645000 ;
      RECT  5.510000 1.755000  5.800000 1.800000 ;
      RECT  5.510000 1.940000  5.800000 1.985000 ;
      RECT  6.090000 0.735000  6.380000 0.780000 ;
      RECT  6.090000 0.920000  6.380000 0.965000 ;
      RECT  6.090000 1.415000  6.380000 1.460000 ;
      RECT  6.090000 1.600000  6.380000 1.645000 ;
      RECT  6.550000 1.075000  6.840000 1.120000 ;
      RECT  6.550000 1.120000 11.450000 1.260000 ;
      RECT  6.550000 1.260000  6.840000 1.305000 ;
      RECT  8.400000 1.415000  8.690000 1.460000 ;
      RECT  8.400000 1.460000 11.910000 1.600000 ;
      RECT  8.400000 1.600000  8.690000 1.645000 ;
      RECT  8.860000 0.735000  9.150000 0.780000 ;
      RECT  8.860000 0.920000  9.150000 0.965000 ;
      RECT  9.020000 1.755000  9.310000 1.800000 ;
      RECT  9.020000 1.800000 10.750000 1.940000 ;
      RECT  9.020000 1.940000  9.310000 1.985000 ;
      RECT 10.460000 1.755000 10.750000 1.800000 ;
      RECT 10.460000 1.940000 10.750000 1.985000 ;
      RECT 11.160000 1.075000 11.450000 1.120000 ;
      RECT 11.160000 1.260000 11.450000 1.305000 ;
      RECT 11.620000 1.415000 11.910000 1.460000 ;
      RECT 11.620000 1.600000 11.910000 1.645000 ;
  END
END sky130_fd_sc_hd__fah_1
END LIBRARY
