# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a41oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 0.995000 4.205000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.405000 1.075000 6.315000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.560000 1.075000 7.955000 1.300000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.075000 9.975000 1.280000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.745000 1.305000 ;
        RECT 0.105000 1.305000 0.325000 1.965000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.575000 2.155000 1.685000 ;
        RECT 0.515000 1.685000 1.685000 1.745000 ;
        RECT 0.515000 1.745000 0.845000 2.085000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 0.635000 4.015000 0.805000 ;
        RECT 1.350000 1.495000 2.155000 1.575000 ;
        RECT 1.350000 1.745000 1.685000 2.085000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.935000 0.805000 2.155000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.090000  0.085000  0.425000 0.465000 ;
        RECT 0.935000  0.085000  1.265000 0.465000 ;
        RECT 1.775000  0.085000  2.105000 0.465000 ;
        RECT 8.405000  0.085000  8.735000 0.465000 ;
        RECT 9.245000  0.085000  9.575000 0.465000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 2.505000 2.255000  3.175000 2.635000 ;
        RECT 3.685000 1.915000  4.015000 2.635000 ;
        RECT 4.620000 1.915000  4.950000 2.635000 ;
        RECT 5.495000 1.915000  6.165000 2.635000 ;
        RECT 6.725000 1.915000  7.055000 2.635000 ;
        RECT 7.565000 1.915000  7.895000 2.635000 ;
        RECT 8.405000 1.915000  8.735000 2.635000 ;
        RECT 9.245000 1.915000  9.575000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 2.255000 2.335000 2.425000 ;
      RECT 2.165000 1.905000 3.515000 2.075000 ;
      RECT 2.165000 2.075000 2.335000 2.255000 ;
      RECT 2.165000 2.425000 2.335000 2.465000 ;
      RECT 2.425000 0.295000 6.115000 0.465000 ;
      RECT 3.345000 1.575000 9.945000 1.745000 ;
      RECT 3.345000 1.745000 3.515000 1.905000 ;
      RECT 3.345000 2.075000 3.515000 2.465000 ;
      RECT 4.185000 1.745000 4.355000 2.425000 ;
      RECT 4.525000 0.635000 7.895000 0.805000 ;
      RECT 5.120000 1.745000 5.290000 2.465000 ;
      RECT 6.305000 0.295000 8.235000 0.465000 ;
      RECT 6.385000 1.745000 6.555000 2.465000 ;
      RECT 7.225000 1.745000 7.395000 2.465000 ;
      RECT 8.065000 0.255000 8.235000 0.295000 ;
      RECT 8.065000 0.465000 8.235000 0.635000 ;
      RECT 8.065000 0.635000 9.915000 0.805000 ;
      RECT 8.065000 1.745000 8.235000 2.465000 ;
      RECT 8.905000 0.255000 9.075000 0.635000 ;
      RECT 8.905000 1.745000 9.075000 2.465000 ;
      RECT 9.745000 0.255000 9.915000 0.635000 ;
      RECT 9.775000 1.745000 9.945000 2.465000 ;
  END
END sky130_fd_sc_hd__a41oi_4
END LIBRARY
