# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__or2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.765000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.835000 2.215000 2.005000 ;
        RECT 1.440000 2.005000 1.770000 2.465000 ;
        RECT 1.520000 0.385000 1.690000 0.655000 ;
        RECT 1.520000 0.655000 2.215000 0.825000 ;
        RECT 1.785000 0.825000 2.215000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.300000 0.085000 ;
        RECT 0.105000  0.085000 0.345000 0.595000 ;
        RECT 1.035000  0.085000 1.350000 0.595000 ;
        RECT 1.860000  0.085000 2.190000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.300000 2.805000 ;
        RECT 1.100000 1.835000 1.270000 2.635000 ;
        RECT 1.940000 2.175000 2.110000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.155000 1.495000 1.615000 1.665000 ;
      RECT 0.155000 1.665000 0.515000 1.840000 ;
      RECT 0.515000 0.255000 0.805000 0.595000 ;
      RECT 0.515000 0.595000 0.695000 1.495000 ;
      RECT 1.445000 0.995000 1.615000 1.495000 ;
  END
END sky130_fd_sc_hd__or2_2
END LIBRARY
