# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.170000 1.075000 7.940000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 1.075000 5.980000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.075000 4.020000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.700000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 2.160000 0.905000 ;
        RECT 0.515000 1.445000 3.885000 1.615000 ;
        RECT 0.515000 1.615000 0.845000 2.465000 ;
        RECT 1.355000 1.615000 1.685000 2.465000 ;
        RECT 1.870000 0.905000 2.160000 1.445000 ;
        RECT 2.715000 1.615000 3.045000 2.125000 ;
        RECT 3.555000 1.615000 3.885000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 2.795000  0.085000  2.965000 0.545000 ;
        RECT 3.635000  0.085000  3.805000 0.545000 ;
        RECT 4.475000  0.085000  4.645000 0.545000 ;
        RECT 5.315000  0.085000  5.485000 0.545000 ;
        RECT 6.675000  0.085000  6.845000 0.545000 ;
        RECT 7.515000  0.085000  7.685000 0.545000 ;
        RECT 8.355000  0.085000  8.525000 0.545000 ;
        RECT 9.195000  0.085000  9.365000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.085000 1.445000  0.345000 2.635000 ;
        RECT 1.015000 1.835000  1.185000 2.635000 ;
        RECT 1.855000 1.835000  2.105000 2.635000 ;
        RECT 8.355000 1.835000  8.525000 2.635000 ;
        RECT 9.195000 1.835000  9.365000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 2.625000 0.465000 ;
      RECT 0.085000 0.465000 0.345000 0.905000 ;
      RECT 2.295000 1.785000 2.545000 2.295000 ;
      RECT 2.295000 2.295000 4.225000 2.465000 ;
      RECT 2.350000 0.465000 2.625000 0.735000 ;
      RECT 2.350000 0.735000 9.865000 0.905000 ;
      RECT 3.135000 0.255000 3.465000 0.735000 ;
      RECT 3.215000 1.785000 3.385000 2.295000 ;
      RECT 3.975000 0.255000 4.305000 0.735000 ;
      RECT 4.055000 1.445000 5.985000 1.615000 ;
      RECT 4.055000 1.615000 4.225000 2.295000 ;
      RECT 4.395000 1.785000 4.645000 2.295000 ;
      RECT 4.395000 2.295000 7.685000 2.465000 ;
      RECT 4.815000 0.255000 5.145000 0.735000 ;
      RECT 4.815000 1.615000 5.145000 2.125000 ;
      RECT 5.315000 1.785000 5.485000 2.295000 ;
      RECT 5.655000 0.255000 5.985000 0.735000 ;
      RECT 5.655000 1.615000 5.985000 2.125000 ;
      RECT 6.175000 0.260000 6.505000 0.735000 ;
      RECT 6.175000 1.445000 9.865000 1.615000 ;
      RECT 6.175000 1.615000 6.505000 2.125000 ;
      RECT 6.675000 1.785000 6.845000 2.295000 ;
      RECT 7.015000 0.260000 7.345000 0.735000 ;
      RECT 7.015000 1.615000 7.345000 2.125000 ;
      RECT 7.515000 1.785000 7.685000 2.295000 ;
      RECT 7.855000 0.260000 8.185000 0.735000 ;
      RECT 7.855000 1.615000 8.185000 2.465000 ;
      RECT 8.695000 0.260000 9.025000 0.735000 ;
      RECT 8.695000 1.615000 9.025000 2.465000 ;
      RECT 9.535000 0.260000 9.865000 0.735000 ;
      RECT 9.535000 1.615000 9.865000 2.465000 ;
  END
END sky130_fd_sc_hd__o41ai_4
END LIBRARY
