# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a32oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.230000 1.075000 1.595000 1.255000 ;
        RECT 1.405000 0.345000 1.705000 0.765000 ;
        RECT 1.405000 0.765000 1.595000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.995000 2.165000 1.325000 ;
        RECT 1.965000 0.415000 2.165000 0.995000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.015000 2.750000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.995000 1.025000 1.425000 ;
        RECT 0.855000 1.425000 1.255000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.575500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 1.165000 0.805000 ;
        RECT 0.515000 0.805000 0.685000 1.785000 ;
        RECT 0.515000 1.785000 0.865000 2.085000 ;
        RECT 0.915000 0.295000 1.165000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.465000 ;
        RECT 2.355000  0.085000 2.695000 0.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 1.555000 2.135000 1.805000 2.635000 ;
        RECT 2.355000 1.495000 2.695000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.835000 0.345000 2.255000 ;
      RECT 0.085000 2.255000 1.345000 2.465000 ;
      RECT 1.095000 1.785000 2.185000 1.955000 ;
      RECT 1.095000 1.955000 1.345000 2.255000 ;
      RECT 2.015000 1.745000 2.185000 1.785000 ;
      RECT 2.015000 1.955000 2.185000 2.465000 ;
  END
END sky130_fd_sc_hd__a32oi_1
END LIBRARY
