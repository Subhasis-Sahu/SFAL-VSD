# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__ha_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.315000 3.585000 1.485000 ;
        RECT 3.360000 1.055000 3.585000 1.315000 ;
        RECT 3.360000 1.485000 3.585000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.850000 1.345000 2.155000 1.655000 ;
        RECT 1.850000 1.655000 3.165000 1.825000 ;
        RECT 1.850000 1.825000 2.155000 2.375000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.315000 4.515000 0.825000 ;
        RECT 4.175000 1.565000 4.515000 2.415000 ;
        RECT 4.330000 0.825000 4.515000 1.565000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.315000 0.425000 0.825000 ;
        RECT 0.090000 0.825000 0.320000 1.565000 ;
        RECT 0.090000 1.565000 0.425000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.595000  0.085000 0.790000 0.885000 ;
        RECT 1.875000  0.085000 2.205000 0.465000 ;
        RECT 3.755000  0.085000 4.005000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.595000 1.515000 0.790000 2.275000 ;
        RECT 0.595000 2.275000 1.260000 2.635000 ;
        RECT 2.450000 2.275000 3.120000 2.635000 ;
        RECT 3.755000 2.125000 4.005000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.490000 1.075000 1.130000 1.245000 ;
      RECT 0.960000 0.345000 1.285000 0.675000 ;
      RECT 0.960000 0.675000 1.130000 1.075000 ;
      RECT 0.960000 1.245000 1.130000 1.935000 ;
      RECT 0.960000 1.935000 1.680000 2.105000 ;
      RECT 1.300000 0.975000 3.170000 1.145000 ;
      RECT 1.300000 1.145000 1.470000 1.325000 ;
      RECT 1.510000 2.105000 1.680000 2.355000 ;
      RECT 1.535000 0.345000 1.705000 0.635000 ;
      RECT 1.535000 0.635000 2.545000 0.805000 ;
      RECT 2.375000 0.345000 2.545000 0.635000 ;
      RECT 3.000000 0.345000 3.170000 0.715000 ;
      RECT 3.000000 0.715000 4.005000 0.885000 ;
      RECT 3.000000 0.885000 3.170000 0.975000 ;
      RECT 3.350000 1.785000 4.005000 1.955000 ;
      RECT 3.350000 1.955000 3.520000 2.355000 ;
      RECT 3.835000 0.885000 4.005000 0.995000 ;
      RECT 3.835000 0.995000 4.160000 1.325000 ;
      RECT 3.835000 1.325000 4.005000 1.785000 ;
  END
END sky130_fd_sc_hd__ha_1
END LIBRARY
