# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__bufbuf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.230000 0.260000 3.560000 0.735000 ;
        RECT 3.230000 0.735000 6.815000 0.905000 ;
        RECT 3.230000 1.445000 6.815000 1.615000 ;
        RECT 3.230000 1.615000 3.560000 2.465000 ;
        RECT 4.070000 0.260000 4.400000 0.735000 ;
        RECT 4.070000 1.615000 4.400000 2.465000 ;
        RECT 4.910000 0.260000 5.240000 0.735000 ;
        RECT 4.910000 1.615000 5.240000 2.465000 ;
        RECT 5.750000 0.260000 6.080000 0.735000 ;
        RECT 5.750000 1.615000 6.080000 2.465000 ;
        RECT 6.435000 0.905000 6.815000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.595000  0.085000 0.765000 0.565000 ;
        RECT 2.050000  0.085000 2.220000 0.565000 ;
        RECT 2.890000  0.085000 3.060000 0.565000 ;
        RECT 3.730000  0.085000 3.900000 0.565000 ;
        RECT 4.570000  0.085000 4.740000 0.565000 ;
        RECT 5.410000  0.085000 5.580000 0.565000 ;
        RECT 6.250000  0.085000 6.420000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.595000 1.785000 0.765000 2.635000 ;
        RECT 2.050000 1.785000 2.220000 2.635000 ;
        RECT 2.890000 1.785000 3.060000 2.635000 ;
        RECT 3.730000 1.835000 3.900000 2.635000 ;
        RECT 4.570000 1.835000 4.740000 2.635000 ;
        RECT 5.410000 1.835000 5.580000 2.635000 ;
        RECT 6.250000 1.835000 6.420000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.260000 0.425000 0.735000 ;
      RECT 0.095000 0.735000 0.780000 0.905000 ;
      RECT 0.095000 1.445000 0.780000 1.615000 ;
      RECT 0.095000 1.615000 0.425000 2.160000 ;
      RECT 0.610000 0.905000 0.780000 0.995000 ;
      RECT 0.610000 0.995000 1.040000 1.325000 ;
      RECT 0.610000 1.325000 0.780000 1.445000 ;
      RECT 1.000000 0.260000 1.380000 0.825000 ;
      RECT 1.000000 1.545000 1.380000 2.465000 ;
      RECT 1.210000 0.825000 1.380000 1.075000 ;
      RECT 1.210000 1.075000 2.720000 1.275000 ;
      RECT 1.210000 1.275000 1.380000 1.545000 ;
      RECT 1.550000 0.260000 1.880000 0.735000 ;
      RECT 1.550000 0.735000 3.060000 0.905000 ;
      RECT 1.550000 1.445000 3.060000 1.615000 ;
      RECT 1.550000 1.615000 1.880000 2.465000 ;
      RECT 2.390000 0.260000 2.720000 0.735000 ;
      RECT 2.390000 1.615000 2.720000 2.465000 ;
      RECT 2.890000 0.905000 3.060000 1.075000 ;
      RECT 2.890000 1.075000 5.360000 1.275000 ;
      RECT 2.890000 1.275000 3.060000 1.445000 ;
  END
END sky130_fd_sc_hd__bufbuf_8
END LIBRARY
