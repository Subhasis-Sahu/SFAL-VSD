# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__or4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 0.995000 3.270000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 2.125000 3.120000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 0.415000 4.055000 0.760000 ;
        RECT 3.780000 1.495000 4.055000 2.465000 ;
        RECT 3.885000 0.760000 4.055000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.140000 0.085000 ;
        RECT 0.655000  0.085000 0.825000 0.825000 ;
        RECT 1.470000  0.085000 1.845000 0.485000 ;
        RECT 2.370000  0.085000 2.700000 0.485000 ;
        RECT 3.210000  0.085000 3.590000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.140000 2.805000 ;
        RECT 0.515000 2.205000 0.845000 2.635000 ;
        RECT 3.290000 1.835000 3.570000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.450000 0.400000 0.825000 ;
      RECT 0.085000 0.825000 0.255000 1.865000 ;
      RECT 0.085000 1.865000 1.915000 2.035000 ;
      RECT 0.085000 2.035000 0.345000 2.455000 ;
      RECT 0.990000 1.525000 1.575000 1.695000 ;
      RECT 1.075000 0.450000 1.245000 0.655000 ;
      RECT 1.075000 0.655000 1.575000 0.825000 ;
      RECT 1.405000 0.825000 1.575000 1.075000 ;
      RECT 1.405000 1.075000 1.830000 1.245000 ;
      RECT 1.405000 1.245000 1.575000 1.525000 ;
      RECT 1.510000 2.205000 2.255000 2.375000 ;
      RECT 1.745000 1.415000 2.395000 1.585000 ;
      RECT 1.745000 1.585000 1.915000 1.865000 ;
      RECT 2.015000 0.305000 2.185000 0.655000 ;
      RECT 2.015000 0.655000 3.610000 0.825000 ;
      RECT 2.085000 1.785000 3.120000 1.955000 ;
      RECT 2.085000 1.955000 2.255000 2.205000 ;
      RECT 2.225000 0.995000 2.395000 1.415000 ;
      RECT 2.870000 0.305000 3.040000 0.655000 ;
      RECT 2.950000 1.495000 3.610000 1.665000 ;
      RECT 2.950000 1.665000 3.120000 1.785000 ;
      RECT 3.440000 0.825000 3.610000 0.995000 ;
      RECT 3.440000 0.995000 3.715000 1.325000 ;
      RECT 3.440000 1.325000 3.610000 1.495000 ;
  END
END sky130_fd_sc_hd__or4bb_1
END LIBRARY
