# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o2111ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 1.075000 5.435000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.075000 4.455000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.200000 1.075000 3.185000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.790000 1.325000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.355000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.302000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.615000 0.935000 0.905000 ;
        RECT 0.605000 0.905000 0.865000 1.495000 ;
        RECT 0.605000 1.495000 4.005000 1.665000 ;
        RECT 0.605000 1.665000 0.865000 2.465000 ;
        RECT 1.535000 1.665000 1.725000 2.465000 ;
        RECT 2.395000 1.665000 2.575000 2.465000 ;
        RECT 3.815000 1.665000 4.005000 2.105000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 3.740000  0.085000 4.070000 0.485000 ;
        RECT 4.600000  0.085000 4.930000 0.480000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.175000 1.525000 0.425000 2.635000 ;
        RECT 1.035000 1.835000 1.365000 2.635000 ;
        RECT 1.895000 1.840000 2.225000 2.635000 ;
        RECT 2.755000 1.835000 3.085000 2.635000 ;
        RECT 4.670000 1.855000 4.930000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.260000 1.300000 0.445000 ;
      RECT 0.175000 0.445000 0.435000 0.865000 ;
      RECT 1.115000 0.445000 1.300000 0.735000 ;
      RECT 1.115000 0.735000 2.275000 0.905000 ;
      RECT 1.470000 0.255000 3.210000 0.445000 ;
      RECT 1.470000 0.445000 1.775000 0.530000 ;
      RECT 1.470000 0.530000 1.760000 0.565000 ;
      RECT 1.925000 0.620000 2.275000 0.735000 ;
      RECT 2.450000 0.655000 5.435000 0.840000 ;
      RECT 2.880000 0.445000 3.210000 0.485000 ;
      RECT 3.310000 1.835000 3.570000 2.275000 ;
      RECT 3.310000 2.275000 4.500000 2.465000 ;
      RECT 3.380000 0.365000 3.570000 0.655000 ;
      RECT 4.240000 0.365000 4.430000 0.650000 ;
      RECT 4.240000 0.650000 5.435000 0.655000 ;
      RECT 4.240000 1.515000 5.360000 1.685000 ;
      RECT 4.240000 1.685000 4.500000 2.275000 ;
      RECT 5.100000 0.365000 5.435000 0.650000 ;
      RECT 5.100000 1.685000 5.360000 2.465000 ;
  END
END sky130_fd_sc_hd__o2111ai_2
END LIBRARY
