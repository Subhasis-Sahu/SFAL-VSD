# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.345000 5.895000 0.745000 ;
        RECT 5.635000 1.670000 5.895000 2.455000 ;
        RECT 5.725000 0.745000 5.895000 1.670000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.345000 4.975000 0.995000 ;
        RECT 4.745000 0.995000 5.075000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.325000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.875000  0.085000 2.205000 0.445000 ;
        RECT 3.755000  0.085000 4.025000 0.610000 ;
        RECT 5.155000  0.085000 5.440000 0.715000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.955000 1.835000 2.245000 2.635000 ;
        RECT 3.930000 2.135000 4.445000 2.635000 ;
        RECT 5.135000 1.915000 5.465000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.795000 0.775000 1.965000 ;
      RECT 0.085000 1.965000 0.345000 2.465000 ;
      RECT 0.170000 0.345000 0.345000 0.635000 ;
      RECT 0.170000 0.635000 0.775000 0.805000 ;
      RECT 0.605000 0.805000 0.775000 1.070000 ;
      RECT 0.605000 1.070000 0.835000 1.400000 ;
      RECT 0.605000 1.400000 0.775000 1.795000 ;
      RECT 1.015000 0.345000 1.185000 1.685000 ;
      RECT 1.015000 1.685000 1.235000 2.465000 ;
      RECT 1.430000 1.495000 2.115000 1.665000 ;
      RECT 1.430000 1.665000 1.785000 2.415000 ;
      RECT 1.510000 0.345000 1.705000 0.615000 ;
      RECT 1.510000 0.615000 2.115000 0.765000 ;
      RECT 1.510000 0.765000 2.335000 0.785000 ;
      RECT 1.945000 0.785000 2.335000 1.095000 ;
      RECT 1.945000 1.095000 2.115000 1.495000 ;
      RECT 2.445000 1.355000 2.835000 1.625000 ;
      RECT 2.445000 1.625000 2.760000 1.685000 ;
      RECT 2.690000 0.765000 3.245000 1.095000 ;
      RECT 2.810000 2.255000 3.625000 2.425000 ;
      RECT 2.815000 0.365000 3.585000 0.535000 ;
      RECT 2.900000 1.785000 3.265000 1.995000 ;
      RECT 3.005000 1.095000 3.245000 1.635000 ;
      RECT 3.005000 1.635000 3.265000 1.785000 ;
      RECT 3.415000 0.535000 3.585000 0.995000 ;
      RECT 3.415000 0.995000 4.175000 1.165000 ;
      RECT 3.455000 1.165000 4.175000 1.325000 ;
      RECT 3.455000 1.325000 3.625000 2.255000 ;
      RECT 3.815000 1.535000 5.465000 1.735000 ;
      RECT 3.815000 1.735000 4.965000 1.865000 ;
      RECT 4.195000 0.295000 4.575000 0.805000 ;
      RECT 4.345000 0.805000 4.575000 1.505000 ;
      RECT 4.345000 1.505000 5.465000 1.535000 ;
      RECT 4.625000 1.865000 4.965000 2.435000 ;
      RECT 5.245000 0.995000 5.555000 1.325000 ;
      RECT 5.245000 1.325000 5.465000 1.505000 ;
    LAYER mcon ;
      RECT 0.605000 1.445000 0.775000 1.615000 ;
      RECT 1.065000 1.785000 1.235000 1.955000 ;
      RECT 2.445000 1.445000 2.615000 1.615000 ;
      RECT 2.925000 1.785000 3.095000 1.955000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.675000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.005000 1.755000 1.295000 1.800000 ;
      RECT 1.005000 1.800000 3.155000 1.940000 ;
      RECT 1.005000 1.940000 1.295000 1.985000 ;
      RECT 2.385000 1.415000 2.675000 1.460000 ;
      RECT 2.385000 1.600000 2.675000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_1
END LIBRARY
