# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a32o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.280000 1.075000 5.075000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335000 1.075000 4.030000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 3.105000 1.295000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.630000 1.075000 6.780000 1.625000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.030000 1.075000 7.710000 1.295000 ;
        RECT 7.030000 1.295000 7.225000 1.635000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.635000 1.605000 0.805000 ;
        RECT 0.120000 0.805000 0.340000 1.495000 ;
        RECT 0.120000 1.495000 1.605000 1.665000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 1.665000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.435000 1.665000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.465000 ;
        RECT 0.935000  0.085000 1.265000 0.465000 ;
        RECT 1.775000  0.085000 2.105000 0.465000 ;
        RECT 2.615000  0.085000 2.945000 0.465000 ;
        RECT 6.975000  0.085000 7.305000 0.465000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.095000 1.915000 0.425000 2.635000 ;
        RECT 0.935000 1.915000 1.265000 2.635000 ;
        RECT 1.775000 1.915000 2.105000 2.635000 ;
        RECT 2.615000 2.255000 2.945000 2.635000 ;
        RECT 3.555000 2.255000 3.885000 2.635000 ;
        RECT 4.395000 2.255000 4.725000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.570000 0.995000 1.970000 1.325000 ;
      RECT 1.800000 1.325000 1.970000 1.495000 ;
      RECT 1.800000 1.495000 5.450000 1.665000 ;
      RECT 2.275000 0.255000 2.445000 0.655000 ;
      RECT 2.275000 0.655000 3.885000 0.825000 ;
      RECT 2.275000 1.915000 5.065000 2.085000 ;
      RECT 2.275000 2.085000 2.445000 2.465000 ;
      RECT 3.135000 0.295000 5.145000 0.465000 ;
      RECT 3.215000 2.085000 3.385000 2.465000 ;
      RECT 4.055000 2.085000 4.225000 2.465000 ;
      RECT 4.395000 0.635000 6.425000 0.805000 ;
      RECT 4.895000 2.085000 5.065000 2.255000 ;
      RECT 4.895000 2.255000 7.725000 2.425000 ;
      RECT 5.280000 0.805000 5.450000 1.495000 ;
      RECT 5.280000 1.665000 5.450000 1.905000 ;
      RECT 5.280000 1.905000 6.200000 1.915000 ;
      RECT 5.280000 1.915000 7.305000 2.075000 ;
      RECT 5.670000 0.295000 6.805000 0.465000 ;
      RECT 6.135000 2.075000 7.305000 2.085000 ;
      RECT 6.635000 0.255000 6.805000 0.295000 ;
      RECT 6.635000 0.465000 6.805000 0.645000 ;
      RECT 6.635000 0.645000 7.645000 0.815000 ;
      RECT 7.475000 0.255000 7.645000 0.645000 ;
      RECT 7.475000 1.755000 7.725000 2.255000 ;
  END
END sky130_fd_sc_hd__a32o_4
END LIBRARY
