# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o32ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.290000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.090000 1.075000 7.260000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.770000 1.075000 5.380000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205000 1.075000 3.540000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.685000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 3.380000 0.905000 ;
        RECT 0.515000 1.495000 5.580000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.085000 ;
        RECT 1.355000 1.665000 1.700000 2.085000 ;
        RECT 1.855000 0.905000 2.035000 1.495000 ;
        RECT 4.410000 1.665000 4.740000 2.085000 ;
        RECT 5.250000 1.665000 5.580000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 3.970000  0.085000  4.140000 0.545000 ;
        RECT 4.810000  0.085000  5.140000 0.545000 ;
        RECT 6.170000  0.085000  6.340000 0.545000 ;
        RECT 7.010000  0.085000  7.180000 0.545000 ;
        RECT 8.370000  0.085000  8.540000 0.545000 ;
        RECT 9.210000  0.085000  9.470000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 2.210000 2.175000  2.540000 2.635000 ;
        RECT 3.050000 2.175000  3.380000 2.635000 ;
        RECT 7.870000 1.835000  8.120000 2.635000 ;
        RECT 8.790000 1.835000  8.960000 2.635000 ;
        RECT 9.630000 1.495000 10.035000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000  3.800000 0.465000 ;
      RECT 0.090000 0.465000  0.345000 0.905000 ;
      RECT 0.090000 1.495000  0.345000 2.255000 ;
      RECT 0.090000 2.255000  2.040000 2.465000 ;
      RECT 1.015000 1.835000  1.185000 2.255000 ;
      RECT 1.870000 1.835000  3.800000 2.005000 ;
      RECT 1.870000 2.005000  2.040000 2.255000 ;
      RECT 2.710000 2.005000  2.880000 2.425000 ;
      RECT 3.550000 0.465000  3.800000 0.735000 ;
      RECT 3.550000 0.735000 10.035000 0.905000 ;
      RECT 3.550000 2.005000  3.800000 2.465000 ;
      RECT 3.990000 1.835000  4.240000 2.255000 ;
      RECT 3.990000 2.255000  7.680000 2.465000 ;
      RECT 4.310000 0.255000  4.640000 0.735000 ;
      RECT 4.910000 1.835000  5.080000 2.255000 ;
      RECT 5.310000 0.255000  5.980000 0.735000 ;
      RECT 5.750000 1.835000  5.920000 2.255000 ;
      RECT 6.090000 1.495000  9.460000 1.665000 ;
      RECT 6.090000 1.665000  6.420000 2.085000 ;
      RECT 6.510000 0.255000  6.840000 0.735000 ;
      RECT 6.590000 1.835000  6.760000 2.255000 ;
      RECT 6.930000 1.665000  7.260000 2.085000 ;
      RECT 7.350000 0.255000  8.040000 0.735000 ;
      RECT 7.430000 1.835000  7.680000 2.255000 ;
      RECT 8.290000 1.665000  8.620000 2.465000 ;
      RECT 8.710000 0.255000  9.040000 0.735000 ;
      RECT 9.130000 1.665000  9.460000 2.465000 ;
      RECT 9.645000 0.255000 10.035000 0.735000 ;
  END
END sky130_fd_sc_hd__o32ai_4
END LIBRARY
