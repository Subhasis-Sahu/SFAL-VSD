# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.795000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.255000 0.255000 9.585000 0.790000 ;
        RECT 9.255000 0.790000 9.615000 0.825000 ;
        RECT 9.255000 1.495000 9.615000 1.530000 ;
        RECT 9.255000 1.530000 9.585000 2.430000 ;
        RECT 9.410000 0.825000 9.615000 0.890000 ;
        RECT 9.410000 1.430000 9.615000 1.495000 ;
        RECT 9.445000 0.890000 9.615000 1.430000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.190000 0.265000 11.440000 0.795000 ;
        RECT 11.190000 1.445000 11.440000 2.325000 ;
        RECT 11.235000 0.795000 11.440000 1.445000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535000 1.035000 4.035000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.255000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.085000 0.785000 3.255000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.960000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  1.975000  0.085000  2.305000 0.445000 ;
        RECT  3.765000  0.085000  3.965000 0.525000 ;
        RECT  5.715000  0.085000  6.085000 0.585000 ;
        RECT  7.740000  0.085000  8.110000 0.615000 ;
        RECT  8.895000  0.085000  9.085000 0.695000 ;
        RECT  9.755000  0.085000  9.985000 0.690000 ;
        RECT 10.690000  0.085000 11.020000 0.805000 ;
        RECT 11.610000  0.085000 11.780000 0.955000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.960000 2.805000 ;
        RECT  0.520000 2.135000  0.850000 2.635000 ;
        RECT  1.880000 2.245000  2.210000 2.635000 ;
        RECT  3.760000 2.165000  3.930000 2.635000 ;
        RECT  5.925000 1.835000  6.095000 2.635000 ;
        RECT  7.805000 2.135000  8.110000 2.635000 ;
        RECT  8.895000 1.625000  9.075000 2.635000 ;
        RECT  9.765000 1.615000  9.935000 2.635000 ;
        RECT 10.715000 1.495000 11.020000 2.635000 ;
        RECT 11.610000 1.395000 11.780000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.175000 0.345000  0.345000 0.635000 ;
      RECT  0.175000 0.635000  0.810000 0.805000 ;
      RECT  0.180000 1.795000  0.845000 1.965000 ;
      RECT  0.180000 1.965000  0.350000 2.465000 ;
      RECT  0.615000 0.805000  0.810000 0.970000 ;
      RECT  0.615000 0.970000  0.845000 1.795000 ;
      RECT  1.015000 0.345000  1.245000 0.715000 ;
      RECT  1.020000 0.715000  1.245000 2.465000 ;
      RECT  1.435000 0.275000  1.805000 0.445000 ;
      RECT  1.435000 0.445000  1.605000 1.860000 ;
      RECT  1.435000 1.860000  3.250000 2.075000 ;
      RECT  1.435000 2.075000  1.710000 2.445000 ;
      RECT  2.120000 0.955000  2.465000 1.125000 ;
      RECT  2.120000 1.125000  2.290000 1.860000 ;
      RECT  2.695000 2.245000  3.590000 2.415000 ;
      RECT  2.820000 0.275000  3.595000 0.445000 ;
      RECT  3.080000 1.355000  3.275000 1.685000 ;
      RECT  3.080000 1.685000  3.250000 1.860000 ;
      RECT  3.420000 1.825000  4.375000 1.995000 ;
      RECT  3.420000 1.995000  3.590000 2.245000 ;
      RECT  3.425000 0.445000  3.595000 0.695000 ;
      RECT  3.425000 0.695000  4.375000 0.865000 ;
      RECT  4.205000 0.365000  4.555000 0.535000 ;
      RECT  4.205000 0.535000  4.375000 0.695000 ;
      RECT  4.205000 0.865000  4.375000 1.825000 ;
      RECT  4.205000 1.995000  4.375000 2.065000 ;
      RECT  4.205000 2.065000  4.485000 2.440000 ;
      RECT  4.545000 0.705000  5.125000 1.035000 ;
      RECT  4.545000 1.035000  4.785000 1.905000 ;
      RECT  4.685000 2.190000  5.755000 2.360000 ;
      RECT  4.725000 0.365000  5.465000 0.535000 ;
      RECT  4.975000 1.655000  5.415000 2.010000 ;
      RECT  5.295000 0.535000  5.465000 1.315000 ;
      RECT  5.295000 1.315000  6.095000 1.485000 ;
      RECT  5.585000 1.485000  6.095000 1.575000 ;
      RECT  5.585000 1.575000  5.755000 2.190000 ;
      RECT  5.635000 0.765000  6.435000 1.065000 ;
      RECT  5.635000 1.065000  5.805000 1.095000 ;
      RECT  5.925000 1.245000  6.095000 1.315000 ;
      RECT  6.265000 0.365000  6.725000 0.535000 ;
      RECT  6.265000 0.535000  6.435000 0.765000 ;
      RECT  6.265000 1.065000  6.435000 2.135000 ;
      RECT  6.265000 2.135000  6.515000 2.465000 ;
      RECT  6.605000 0.705000  7.155000 1.035000 ;
      RECT  6.605000 1.245000  6.795000 1.965000 ;
      RECT  6.740000 2.165000  7.625000 2.335000 ;
      RECT  6.955000 0.365000  7.495000 0.535000 ;
      RECT  6.965000 1.035000  7.155000 1.575000 ;
      RECT  6.965000 1.575000  7.285000 1.905000 ;
      RECT  7.325000 0.535000  7.495000 0.995000 ;
      RECT  7.325000 0.995000  8.370000 1.325000 ;
      RECT  7.325000 1.325000  7.625000 1.405000 ;
      RECT  7.455000 1.405000  7.625000 2.165000 ;
      RECT  7.795000 1.575000  8.725000 1.905000 ;
      RECT  8.360000 0.300000  8.725000 0.825000 ;
      RECT  8.395000 1.905000  8.725000 2.455000 ;
      RECT  8.540000 0.825000  8.725000 0.995000 ;
      RECT  8.540000 0.995000  9.275000 1.325000 ;
      RECT  8.540000 1.325000  8.725000 1.575000 ;
      RECT 10.205000 0.345000 10.455000 0.995000 ;
      RECT 10.205000 0.995000 11.065000 1.325000 ;
      RECT 10.205000 1.325000 10.535000 2.425000 ;
    LAYER mcon ;
      RECT 0.645000 1.785000 0.815000 1.955000 ;
      RECT 1.050000 0.765000 1.220000 0.935000 ;
      RECT 4.745000 0.765000 4.915000 0.935000 ;
      RECT 5.205000 1.785000 5.375000 1.955000 ;
      RECT 6.625000 1.785000 6.795000 1.955000 ;
      RECT 6.640000 0.765000 6.810000 0.935000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 6.855000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 0.990000 0.735000 1.280000 0.780000 ;
      RECT 0.990000 0.780000 6.870000 0.920000 ;
      RECT 0.990000 0.920000 1.280000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.565000 1.755000 6.855000 1.800000 ;
      RECT 6.565000 1.940000 6.855000 1.985000 ;
      RECT 6.580000 0.735000 6.870000 0.780000 ;
      RECT 6.580000 0.920000 6.870000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxbp_2
END LIBRARY
