# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__bufbuf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  5.235000 0.255000  5.485000 0.260000 ;
        RECT  5.235000 0.260000  5.565000 0.735000 ;
        RECT  5.235000 0.735000 11.875000 0.905000 ;
        RECT  5.235000 1.445000 11.875000 1.615000 ;
        RECT  5.235000 1.615000  5.565000 2.465000 ;
        RECT  6.075000 0.260000  6.405000 0.735000 ;
        RECT  6.075000 1.615000  6.405000 2.465000 ;
        RECT  6.155000 0.255000  6.325000 0.260000 ;
        RECT  6.915000 0.260000  7.245000 0.735000 ;
        RECT  6.915000 1.615000  7.245000 2.465000 ;
        RECT  6.995000 0.255000  7.165000 0.260000 ;
        RECT  7.755000 0.260000  8.085000 0.735000 ;
        RECT  7.755000 1.615000  8.085000 2.465000 ;
        RECT  8.595000 0.260000  8.925000 0.735000 ;
        RECT  8.595000 1.615000  8.925000 2.465000 ;
        RECT  9.435000 0.260000  9.765000 0.735000 ;
        RECT  9.435000 1.615000  9.765000 2.465000 ;
        RECT 10.275000 0.260000 10.605000 0.735000 ;
        RECT 10.275000 1.615000 10.605000 2.465000 ;
        RECT 11.115000 0.260000 11.445000 0.735000 ;
        RECT 11.115000 1.615000 11.445000 2.465000 ;
        RECT 11.620000 0.905000 11.875000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.960000 0.085000 ;
        RECT  0.175000  0.085000  0.345000 0.905000 ;
        RECT  1.535000  0.085000  1.705000 0.565000 ;
        RECT  2.375000  0.085000  2.545000 0.565000 ;
        RECT  3.215000  0.085000  3.385000 0.565000 ;
        RECT  4.055000  0.085000  4.225000 0.565000 ;
        RECT  4.895000  0.085000  5.065000 0.565000 ;
        RECT  5.735000  0.085000  5.905000 0.565000 ;
        RECT  6.575000  0.085000  6.745000 0.565000 ;
        RECT  7.415000  0.085000  7.585000 0.565000 ;
        RECT  8.255000  0.085000  8.425000 0.565000 ;
        RECT  9.095000  0.085000  9.265000 0.565000 ;
        RECT  9.935000  0.085000 10.105000 0.565000 ;
        RECT 10.775000  0.085000 10.945000 0.565000 ;
        RECT 11.615000  0.085000 11.785000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.960000 2.805000 ;
        RECT  0.175000 1.445000  0.345000 2.635000 ;
        RECT  1.535000 1.785000  1.705000 2.635000 ;
        RECT  2.375000 1.785000  2.545000 2.635000 ;
        RECT  3.215000 1.835000  3.385000 2.635000 ;
        RECT  4.055000 1.835000  4.225000 2.635000 ;
        RECT  4.895000 1.835000  5.065000 2.635000 ;
        RECT  5.735000 1.835000  5.905000 2.635000 ;
        RECT  6.575000 1.835000  6.745000 2.635000 ;
        RECT  7.415000 1.835000  7.585000 2.635000 ;
        RECT  8.255000 1.835000  8.425000 2.635000 ;
        RECT  9.095000 1.835000  9.265000 2.635000 ;
        RECT  9.935000 1.835000 10.105000 2.635000 ;
        RECT 10.775000 1.835000 10.945000 2.635000 ;
        RECT 11.615000 1.835000 11.785000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 0.260000  0.845000 0.905000 ;
      RECT 0.515000 1.445000  0.845000 2.465000 ;
      RECT 0.610000 0.905000  0.845000 1.075000 ;
      RECT 0.610000 1.075000  2.205000 1.275000 ;
      RECT 0.610000 1.275000  0.845000 1.445000 ;
      RECT 1.035000 0.260000  1.365000 0.735000 ;
      RECT 1.035000 0.735000  2.545000 0.905000 ;
      RECT 1.035000 1.445000  2.545000 1.615000 ;
      RECT 1.035000 1.615000  1.365000 2.465000 ;
      RECT 1.875000 0.260000  2.205000 0.735000 ;
      RECT 1.875000 1.615000  2.205000 2.465000 ;
      RECT 2.375000 0.905000  2.545000 1.075000 ;
      RECT 2.375000 1.075000  4.685000 1.275000 ;
      RECT 2.375000 1.275000  2.545000 1.445000 ;
      RECT 2.715000 0.260000  3.045000 0.735000 ;
      RECT 2.715000 0.735000  5.065000 0.905000 ;
      RECT 2.715000 1.445000  5.065000 1.615000 ;
      RECT 2.715000 1.615000  3.045000 2.465000 ;
      RECT 3.555000 0.260000  3.885000 0.735000 ;
      RECT 3.555000 1.615000  3.885000 2.465000 ;
      RECT 4.395000 0.260000  4.725000 0.735000 ;
      RECT 4.395000 1.615000  4.725000 2.465000 ;
      RECT 4.890000 0.905000  5.065000 1.075000 ;
      RECT 4.890000 1.075000 11.450000 1.275000 ;
      RECT 4.890000 1.275000  5.065000 1.445000 ;
  END
END sky130_fd_sc_hd__bufbuf_16
END LIBRARY
