# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__fa_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.080000 0.995000 2.680000 1.275000 ;
        RECT 2.080000 1.275000 2.340000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.610000 1.030000 4.000000 1.360000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.645000 0.955000 6.005000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.030000 0.995000 7.885000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.390000 1.075000 2.680000 1.120000 ;
        RECT 2.390000 1.120000 7.300000 1.260000 ;
        RECT 2.390000 1.260000 2.680000 1.305000 ;
        RECT 3.770000 1.075000 4.060000 1.120000 ;
        RECT 3.770000 1.260000 4.060000 1.305000 ;
        RECT 5.630000 1.075000 5.920000 1.120000 ;
        RECT 5.630000 1.260000 5.920000 1.305000 ;
        RECT 7.010000 1.075000 7.300000 1.120000 ;
        RECT 7.010000 1.260000 7.300000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 1.445000 3.080000 1.690000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.580000 1.435000 4.995000 1.745000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.075000 1.445000 7.760000 1.735000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.850000 1.415000 3.140000 1.460000 ;
        RECT 2.850000 1.460000 7.760000 1.600000 ;
        RECT 2.850000 1.600000 3.140000 1.645000 ;
        RECT 4.710000 1.415000 5.000000 1.460000 ;
        RECT 4.710000 1.600000 5.000000 1.645000 ;
        RECT 7.470000 1.415000 7.760000 1.460000 ;
        RECT 7.470000 1.600000 7.760000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.105000 3.420000 1.275000 ;
        RECT 3.250000 1.275000 3.420000 1.570000 ;
        RECT 3.250000 1.570000 4.340000 1.740000 ;
        RECT 4.170000 0.965000 5.390000 1.250000 ;
        RECT 4.170000 1.250000 4.340000 1.570000 ;
        RECT 5.220000 1.250000 5.390000 1.435000 ;
        RECT 5.220000 1.435000 5.580000 1.515000 ;
        RECT 5.220000 1.515000 6.845000 1.685000 ;
        RECT 6.595000 1.355000 6.845000 1.515000 ;
        RECT 6.595000 1.685000 6.845000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.735000 1.525000 0.905000 ;
        RECT 0.085000 0.905000 0.435000 1.415000 ;
        RECT 0.085000 1.415000 1.570000 1.585000 ;
        RECT 0.515000 0.255000 0.845000 0.735000 ;
        RECT 0.515000 1.585000 0.845000 2.445000 ;
        RECT 1.355000 0.315000 1.685000 0.485000 ;
        RECT 1.355000 0.485000 1.525000 0.735000 ;
        RECT 1.400000 1.585000 1.570000 1.780000 ;
        RECT 1.400000 1.780000 1.645000 1.950000 ;
        RECT 1.435000 1.950000 1.645000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.943000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.320000 0.255000  8.650000 0.485000 ;
        RECT 8.320000 1.795000  8.570000 1.965000 ;
        RECT 8.320000 1.965000  8.490000 2.465000 ;
        RECT 8.400000 0.485000  8.650000 0.735000 ;
        RECT 8.400000 0.735000 10.035000 0.905000 ;
        RECT 8.400000 1.415000 10.035000 1.585000 ;
        RECT 8.400000 1.585000  8.570000 1.795000 ;
        RECT 9.160000 0.270000  9.490000 0.735000 ;
        RECT 9.160000 1.585000  9.490000 2.425000 ;
        RECT 9.700000 0.905000 10.035000 1.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.175000  0.085000  0.345000 0.565000 ;
        RECT 1.015000  0.085000  1.185000 0.565000 ;
        RECT 1.855000  0.085000  2.185000 0.465000 ;
        RECT 3.680000  0.085000  4.010000 0.445000 ;
        RECT 4.620000  0.085000  4.950000 0.490000 ;
        RECT 5.460000  0.085000  5.790000 0.445000 ;
        RECT 7.705000  0.085000  8.035000 0.445000 ;
        RECT 8.820000  0.085000  8.990000 0.565000 ;
        RECT 9.660000  0.085000  9.830000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.175000 1.795000  0.345000 2.635000 ;
        RECT 1.015000 1.795000  1.185000 2.635000 ;
        RECT 1.815000 2.275000  2.145000 2.635000 ;
        RECT 3.680000 2.275000  4.010000 2.635000 ;
        RECT 4.620000 1.915000  4.950000 2.635000 ;
        RECT 5.460000 2.275000  5.790000 2.635000 ;
        RECT 7.815000 2.275000  8.145000 2.635000 ;
        RECT 8.740000 1.795000  8.910000 2.635000 ;
        RECT 9.660000 1.795000  9.830000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.605000 1.075000 1.910000 1.245000 ;
      RECT 1.740000 0.655000 3.090000 0.825000 ;
      RECT 1.740000 0.825000 1.910000 1.075000 ;
      RECT 1.740000 1.245000 1.910000 1.430000 ;
      RECT 1.740000 1.430000 1.945000 1.495000 ;
      RECT 1.740000 1.495000 2.310000 1.600000 ;
      RECT 1.775000 1.600000 2.310000 1.665000 ;
      RECT 2.140000 1.665000 2.310000 1.910000 ;
      RECT 2.140000 1.910000 3.170000 2.080000 ;
      RECT 2.370000 0.255000 3.090000 0.655000 ;
      RECT 2.735000 2.080000 3.170000 2.465000 ;
      RECT 2.850000 0.825000 3.090000 0.935000 ;
      RECT 3.340000 0.255000 3.510000 0.615000 ;
      RECT 3.340000 0.615000 4.350000 0.785000 ;
      RECT 3.340000 1.935000 4.415000 2.105000 ;
      RECT 3.340000 2.105000 3.510000 2.465000 ;
      RECT 4.180000 0.255000 4.350000 0.615000 ;
      RECT 4.180000 2.105000 4.415000 2.465000 ;
      RECT 5.120000 0.255000 5.290000 0.615000 ;
      RECT 5.120000 0.615000 6.130000 0.785000 ;
      RECT 5.120000 1.935000 6.130000 2.105000 ;
      RECT 5.120000 2.105000 5.290000 2.465000 ;
      RECT 5.960000 0.255000 6.130000 0.615000 ;
      RECT 5.960000 2.105000 6.130000 2.465000 ;
      RECT 6.175000 0.955000 6.860000 1.125000 ;
      RECT 6.345000 0.765000 6.860000 0.955000 ;
      RECT 6.410000 2.125000 7.610000 2.465000 ;
      RECT 6.465000 0.255000 7.475000 0.505000 ;
      RECT 6.465000 0.505000 6.635000 0.595000 ;
      RECT 7.305000 0.505000 7.475000 0.655000 ;
      RECT 7.305000 0.655000 8.225000 0.825000 ;
      RECT 7.440000 1.935000 8.105000 2.105000 ;
      RECT 7.440000 2.105000 7.610000 2.125000 ;
      RECT 7.935000 1.470000 8.225000 1.640000 ;
      RECT 7.935000 1.640000 8.105000 1.935000 ;
      RECT 8.055000 0.825000 8.225000 1.075000 ;
      RECT 8.055000 1.075000 9.445000 1.245000 ;
      RECT 8.055000 1.245000 8.225000 1.470000 ;
    LAYER mcon ;
      RECT 2.910000 0.765000 3.080000 0.935000 ;
      RECT 6.610000 0.765000 6.780000 0.935000 ;
    LAYER met1 ;
      RECT 2.850000 0.735000 3.140000 0.780000 ;
      RECT 2.850000 0.780000 6.840000 0.920000 ;
      RECT 2.850000 0.920000 3.140000 0.965000 ;
      RECT 6.550000 0.735000 6.840000 0.780000 ;
      RECT 6.550000 0.920000 6.840000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_4
END LIBRARY
