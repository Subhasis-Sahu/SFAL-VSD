# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__bufinv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.505000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 0.260000 3.045000 0.735000 ;
        RECT 2.715000 0.735000 6.355000 0.905000 ;
        RECT 2.715000 1.445000 6.355000 1.615000 ;
        RECT 2.715000 1.615000 3.045000 2.465000 ;
        RECT 3.555000 0.260000 3.885000 0.735000 ;
        RECT 3.555000 1.615000 3.885000 2.465000 ;
        RECT 4.395000 0.260000 4.725000 0.735000 ;
        RECT 4.395000 1.615000 4.725000 2.465000 ;
        RECT 5.235000 0.260000 5.565000 0.735000 ;
        RECT 5.235000 1.615000 5.565000 2.465000 ;
        RECT 5.970000 0.905000 6.355000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.175000  0.085000 0.345000 0.905000 ;
        RECT 1.535000  0.085000 1.705000 0.565000 ;
        RECT 2.375000  0.085000 2.545000 0.565000 ;
        RECT 3.215000  0.085000 3.385000 0.565000 ;
        RECT 4.055000  0.085000 4.225000 0.565000 ;
        RECT 4.895000  0.085000 5.065000 0.565000 ;
        RECT 5.735000  0.085000 5.905000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.175000 1.445000 0.345000 2.635000 ;
        RECT 1.535000 1.785000 1.705000 2.635000 ;
        RECT 2.375000 1.785000 2.545000 2.635000 ;
        RECT 3.215000 1.835000 3.385000 2.635000 ;
        RECT 4.055000 1.835000 4.225000 2.635000 ;
        RECT 4.895000 1.835000 5.065000 2.635000 ;
        RECT 5.735000 1.835000 5.905000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 0.260000 0.845000 0.905000 ;
      RECT 0.515000 1.545000 0.845000 2.465000 ;
      RECT 0.675000 0.905000 0.845000 1.075000 ;
      RECT 0.675000 1.075000 2.205000 1.275000 ;
      RECT 0.675000 1.275000 0.845000 1.545000 ;
      RECT 1.035000 0.260000 1.365000 0.735000 ;
      RECT 1.035000 0.735000 2.545000 0.905000 ;
      RECT 1.035000 1.445000 2.545000 1.615000 ;
      RECT 1.035000 1.615000 1.365000 2.465000 ;
      RECT 1.875000 0.260000 2.205000 0.735000 ;
      RECT 1.875000 1.615000 2.205000 2.465000 ;
      RECT 2.375000 0.905000 2.545000 1.075000 ;
      RECT 2.375000 1.075000 5.760000 1.275000 ;
      RECT 2.375000 1.275000 2.545000 1.445000 ;
  END
END sky130_fd_sc_hd__bufinv_8
END LIBRARY
