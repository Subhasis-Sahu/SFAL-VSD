# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nand4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.170000 0.890000 1.340000 ;
        RECT 0.610000 1.070000 0.890000 1.170000 ;
        RECT 0.610000 1.340000 0.890000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.070000 0.330000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.615000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.075000 5.875000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085000 0.655000 2.415000 1.445000 ;
        RECT 2.085000 1.445000 5.455000 1.665000 ;
        RECT 2.085000 1.665000 2.335000 2.465000 ;
        RECT 2.925000 1.665000 3.255000 2.465000 ;
        RECT 3.245000 1.075000 3.550000 1.445000 ;
        RECT 4.285000 1.665000 4.615000 2.465000 ;
        RECT 5.125000 1.665000 5.455000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.515000  0.085000 0.765000 0.545000 ;
        RECT 5.205000  0.085000 5.375000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.540000 2.195000 0.765000 2.635000 ;
        RECT 1.745000 1.495000 1.915000 2.635000 ;
        RECT 2.505000 1.835000 2.755000 2.635000 ;
        RECT 3.425000 1.835000 4.115000 2.635000 ;
        RECT 4.785000 1.835000 4.955000 2.635000 ;
        RECT 5.625000 1.445000 5.895000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.345000 0.730000 ;
      RECT 0.085000 0.730000 1.230000 0.900000 ;
      RECT 0.085000 1.785000 1.230000 1.980000 ;
      RECT 0.085000 1.980000 0.370000 2.440000 ;
      RECT 0.935000 0.255000 1.575000 0.560000 ;
      RECT 0.935000 2.150000 1.575000 2.465000 ;
      RECT 1.060000 0.900000 1.230000 1.785000 ;
      RECT 1.400000 0.560000 1.575000 0.715000 ;
      RECT 1.400000 0.715000 1.580000 1.410000 ;
      RECT 1.400000 1.410000 1.575000 2.150000 ;
      RECT 1.745000 0.255000 3.675000 0.485000 ;
      RECT 1.745000 0.485000 1.915000 0.585000 ;
      RECT 2.745000 1.075000 3.075000 1.275000 ;
      RECT 2.925000 0.655000 4.615000 0.905000 ;
      RECT 3.865000 0.255000 5.035000 0.485000 ;
      RECT 4.785000 0.485000 5.035000 0.735000 ;
      RECT 4.785000 0.735000 5.895000 0.905000 ;
      RECT 5.545000 0.255000 5.895000 0.735000 ;
    LAYER mcon ;
      RECT 1.060000 1.105000 1.230000 1.275000 ;
      RECT 2.905000 1.105000 3.075000 1.275000 ;
    LAYER met1 ;
      RECT 1.000000 1.075000 3.135000 1.305000 ;
  END
END sky130_fd_sc_hd__nand4bb_2
END LIBRARY
