# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a2bb2oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 1.075000 7.320000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595000 1.075000 9.045000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.555000 1.285000 ;
        RECT 1.385000 1.285000 1.555000 1.445000 ;
        RECT 1.385000 1.445000 3.575000 1.615000 ;
        RECT 3.245000 1.075000 3.575000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725000 1.075000 3.075000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 0.645000 2.995000 0.725000 ;
        RECT 1.775000 0.725000 5.045000 0.905000 ;
        RECT 3.745000 0.905000 3.915000 1.415000 ;
        RECT 3.745000 1.415000 4.965000 1.615000 ;
        RECT 3.875000 0.275000 4.205000 0.725000 ;
        RECT 3.915000 1.615000 4.165000 2.125000 ;
        RECT 4.715000 0.275000 5.045000 0.725000 ;
        RECT 4.745000 1.615000 4.965000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.175000  0.085000 0.345000 0.895000 ;
        RECT 1.015000  0.085000 1.185000 0.555000 ;
        RECT 3.535000  0.085000 3.705000 0.555000 ;
        RECT 4.375000  0.085000 4.545000 0.555000 ;
        RECT 5.215000  0.085000 5.905000 0.555000 ;
        RECT 6.575000  0.085000 6.745000 0.555000 ;
        RECT 7.415000  0.085000 7.585000 0.555000 ;
        RECT 8.255000  0.085000 8.425000 0.555000 ;
        RECT 9.095000  0.085000 9.265000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.595000 1.795000 0.805000 2.635000 ;
        RECT 1.395000 2.135000 1.645000 2.635000 ;
        RECT 2.235000 2.135000 2.485000 2.635000 ;
        RECT 3.075000 2.135000 3.325000 2.635000 ;
        RECT 6.155000 1.795000 6.365000 2.635000 ;
        RECT 6.955000 1.795000 7.205000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.455000 1.215000 1.625000 ;
      RECT 0.085000 1.625000 0.425000 2.465000 ;
      RECT 0.515000 0.255000 0.845000 0.725000 ;
      RECT 0.515000 0.725000 1.605000 0.905000 ;
      RECT 0.975000 1.625000 1.215000 1.795000 ;
      RECT 0.975000 1.795000 3.745000 1.965000 ;
      RECT 0.975000 1.965000 1.215000 2.465000 ;
      RECT 1.355000 0.255000 3.365000 0.475000 ;
      RECT 1.355000 0.475000 1.605000 0.725000 ;
      RECT 1.815000 1.965000 2.065000 2.465000 ;
      RECT 2.655000 1.965000 2.905000 2.465000 ;
      RECT 3.495000 1.965000 3.745000 2.295000 ;
      RECT 3.495000 2.295000 5.465000 2.465000 ;
      RECT 4.085000 1.075000 5.725000 1.245000 ;
      RECT 4.335000 1.795000 4.575000 2.295000 ;
      RECT 5.135000 1.455000 5.465000 2.295000 ;
      RECT 5.555000 0.735000 9.575000 0.905000 ;
      RECT 5.555000 0.905000 5.725000 1.075000 ;
      RECT 5.655000 1.455000 7.625000 1.625000 ;
      RECT 5.655000 1.625000 5.985000 2.465000 ;
      RECT 6.075000 0.255000 6.405000 0.725000 ;
      RECT 6.075000 0.725000 8.925000 0.735000 ;
      RECT 6.540000 1.625000 6.780000 2.465000 ;
      RECT 6.915000 0.255000 7.245000 0.725000 ;
      RECT 7.375000 1.625000 7.625000 2.295000 ;
      RECT 7.375000 2.295000 9.310000 2.465000 ;
      RECT 7.755000 0.255000 8.085000 0.725000 ;
      RECT 7.795000 1.455000 9.575000 1.625000 ;
      RECT 7.795000 1.625000 8.045000 2.125000 ;
      RECT 8.215000 1.795000 8.465000 2.295000 ;
      RECT 8.595000 0.255000 8.925000 0.725000 ;
      RECT 8.635000 1.625000 8.885000 2.125000 ;
      RECT 9.060000 1.795000 9.310000 2.295000 ;
      RECT 9.215000 0.905000 9.575000 1.455000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_4
END LIBRARY
