VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pfd_lay
  CLASS BLOCK ;
  FOREIGN pfd_lay ;
  ORIGIN -3.250 15.880 ;
  SIZE 34.000 BY 22.490 ;
  PIN f_clk_in
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 6.950 2.900 7.280 2.915 ;
        RECT 5.950 2.700 7.280 2.900 ;
        RECT 6.950 2.675 7.280 2.700 ;
      LAYER met1 ;
        RECT 4.250 2.900 5.250 3.380 ;
        RECT 5.920 2.900 6.180 2.960 ;
        RECT 4.250 2.700 6.180 2.900 ;
        RECT 4.250 2.380 5.250 2.700 ;
        RECT 5.920 2.640 6.180 2.700 ;
    END
  END f_clk_in
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.440 2.905 27.520 4.510 ;
      LAYER li1 ;
        RECT 6.630 4.235 8.010 4.405 ;
        RECT 10.310 4.235 11.690 4.405 ;
        RECT 14.450 4.235 15.830 4.405 ;
        RECT 17.670 4.235 19.050 4.405 ;
        RECT 21.350 4.235 23.190 4.405 ;
        RECT 25.490 4.235 27.330 4.405 ;
        RECT 6.970 3.095 7.180 4.235 ;
        RECT 10.395 3.095 10.675 4.235 ;
        RECT 11.345 3.095 11.605 4.235 ;
        RECT 14.790 3.095 15.000 4.235 ;
        RECT 18.010 3.095 18.220 4.235 ;
        RECT 21.440 3.095 21.695 4.235 ;
        RECT 22.365 3.435 22.595 4.235 ;
        RECT 25.830 3.095 26.040 4.235 ;
        RECT 26.955 3.070 27.245 4.235 ;
      LAYER met1 ;
        RECT 16.560 5.240 17.560 6.100 ;
        RECT 6.900 4.760 27.040 5.240 ;
        RECT 6.900 4.560 27.600 4.760 ;
        RECT 6.630 4.420 27.600 4.560 ;
        RECT 6.630 4.080 8.010 4.420 ;
        RECT 10.310 4.080 11.690 4.420 ;
        RECT 14.450 4.080 15.830 4.420 ;
        RECT 17.670 4.080 19.050 4.420 ;
        RECT 21.350 4.080 23.190 4.420 ;
        RECT 25.490 4.080 27.330 4.420 ;
    END
    PORT
      LAYER nwell ;
        RECT 19.900 -2.905 23.660 -1.300 ;
      LAYER li1 ;
        RECT 20.090 -1.575 22.390 -1.405 ;
        RECT 23.010 -1.575 23.470 -1.405 ;
        RECT 20.175 -2.715 20.435 -1.575 ;
        RECT 21.105 -2.375 21.275 -1.575 ;
        RECT 22.005 -2.375 22.285 -1.575 ;
        RECT 23.095 -2.740 23.385 -1.575 ;
      LAYER met1 ;
        RECT 20.800 -1.250 21.800 -0.500 ;
        RECT 20.090 -1.730 23.470 -1.250 ;
        RECT 22.250 -1.750 23.220 -1.730 ;
    END
    PORT
      LAYER nwell ;
        RECT 10.580 -13.075 14.550 -13.015 ;
        RECT 10.580 -13.145 15.570 -13.075 ;
        RECT 10.580 -14.620 16.240 -13.145 ;
        RECT 13.810 -14.680 16.240 -14.620 ;
        RECT 15.400 -14.750 16.240 -14.680 ;
      LAYER li1 ;
        RECT 10.855 -14.345 11.115 -13.205 ;
        RECT 11.785 -14.345 12.065 -13.205 ;
        RECT 10.770 -14.515 12.150 -14.345 ;
        RECT 14.085 -14.405 14.345 -13.265 ;
        RECT 15.015 -14.405 15.295 -13.265 ;
        RECT 14.000 -14.575 15.380 -14.405 ;
        RECT 15.675 -14.475 15.965 -13.310 ;
        RECT 15.590 -14.645 16.050 -14.475 ;
      LAYER met1 ;
        RECT 10.770 -14.620 12.150 -14.190 ;
        RECT 14.000 -14.620 15.380 -14.250 ;
        RECT 15.590 -14.620 16.050 -14.320 ;
        RECT 10.580 -14.800 16.050 -14.620 ;
        RECT 10.580 -14.960 15.640 -14.800 ;
        RECT 13.340 -15.880 14.340 -14.960 ;
    END
    PORT
      LAYER nwell ;
        RECT 27.890 -8.410 28.730 -8.400 ;
        RECT 7.360 -10.005 28.730 -8.410 ;
        RECT 7.360 -10.015 27.980 -10.005 ;
      LAYER li1 ;
        RECT 7.550 -8.685 8.930 -8.515 ;
        RECT 11.230 -8.685 12.610 -8.515 ;
        RECT 15.370 -8.685 16.750 -8.515 ;
        RECT 18.590 -8.685 19.970 -8.515 ;
        RECT 22.270 -8.685 24.110 -8.515 ;
        RECT 26.410 -8.685 27.790 -8.515 ;
        RECT 28.080 -8.675 28.540 -8.505 ;
        RECT 7.890 -9.825 8.100 -8.685 ;
        RECT 11.315 -9.825 11.595 -8.685 ;
        RECT 12.265 -9.825 12.525 -8.685 ;
        RECT 15.710 -9.825 15.920 -8.685 ;
        RECT 18.930 -9.825 19.140 -8.685 ;
        RECT 22.360 -9.825 22.615 -8.685 ;
        RECT 23.285 -9.485 23.515 -8.685 ;
        RECT 26.750 -9.825 26.960 -8.685 ;
        RECT 28.165 -9.840 28.455 -8.675 ;
      LAYER met1 ;
        RECT 17.940 -8.025 18.940 -7.160 ;
        RECT 7.830 -8.160 27.970 -8.025 ;
        RECT 7.830 -8.350 28.520 -8.160 ;
        RECT 7.830 -8.360 28.540 -8.350 ;
        RECT 7.550 -8.830 28.540 -8.360 ;
        RECT 7.550 -8.840 28.150 -8.830 ;
        RECT 7.830 -8.845 28.150 -8.840 ;
        RECT 27.900 -8.850 28.150 -8.845 ;
    END
    PORT
      LAYER nwell ;
        RECT 13.120 -0.655 14.880 -0.605 ;
        RECT 9.270 -0.660 11.300 -0.655 ;
        RECT 12.570 -0.660 14.880 -0.655 ;
        RECT 9.270 -0.675 14.880 -0.660 ;
        RECT 8.630 -2.210 14.880 -0.675 ;
        RECT 8.630 -2.260 13.580 -2.210 ;
        RECT 8.630 -2.280 9.470 -2.260 ;
      LAYER li1 ;
        RECT 8.905 -2.005 9.195 -0.840 ;
        RECT 9.545 -1.985 9.825 -0.845 ;
        RECT 10.495 -1.985 10.755 -0.845 ;
        RECT 13.395 -1.935 13.675 -0.795 ;
        RECT 14.345 -1.935 14.605 -0.795 ;
        RECT 8.820 -2.175 9.280 -2.005 ;
        RECT 9.460 -2.155 10.840 -1.985 ;
        RECT 13.310 -2.105 14.690 -1.935 ;
      LAYER met1 ;
        RECT 8.820 -2.040 9.280 -1.850 ;
        RECT 9.460 -2.040 10.840 -1.830 ;
        RECT 13.310 -2.040 14.690 -1.780 ;
        RECT 8.820 -2.330 15.180 -2.040 ;
        RECT 9.200 -2.720 15.180 -2.330 ;
        RECT 12.420 -3.400 13.420 -2.720 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 26.885 1.790 27.315 2.575 ;
        RECT 8.835 -0.345 9.265 0.440 ;
      LAYER li1 ;
        RECT 6.950 1.685 7.180 2.505 ;
        RECT 10.395 1.685 10.705 2.485 ;
        RECT 14.770 1.685 15.000 2.505 ;
        RECT 17.990 1.685 18.220 2.505 ;
        RECT 21.440 1.685 21.695 2.175 ;
        RECT 25.810 1.685 26.040 2.505 ;
        RECT 26.955 1.685 27.245 2.410 ;
        RECT 6.630 1.515 8.010 1.685 ;
        RECT 10.310 1.515 11.690 1.685 ;
        RECT 14.450 1.515 15.830 1.685 ;
        RECT 17.670 1.515 19.050 1.685 ;
        RECT 21.350 1.515 23.190 1.685 ;
        RECT 25.490 1.515 27.330 1.685 ;
        RECT 8.820 0.545 9.280 0.715 ;
        RECT 9.460 0.565 10.840 0.735 ;
        RECT 13.310 0.615 14.690 0.785 ;
        RECT 8.905 -0.180 9.195 0.545 ;
        RECT 9.545 -0.235 9.855 0.565 ;
        RECT 13.395 -0.185 13.705 0.615 ;
      LAYER met1 ;
        RECT 6.630 1.500 8.010 1.840 ;
        RECT 10.310 1.500 11.690 1.840 ;
        RECT 14.450 1.500 15.830 1.840 ;
        RECT 17.670 1.500 19.050 1.840 ;
        RECT 21.350 1.500 23.190 1.840 ;
        RECT 25.490 1.500 27.330 1.840 ;
        RECT 6.630 1.360 27.330 1.500 ;
        RECT 6.900 1.020 27.600 1.360 ;
        RECT 6.900 0.680 27.040 1.020 ;
        RECT 8.820 0.390 9.280 0.680 ;
        RECT 9.460 0.410 10.840 0.680 ;
        RECT 13.310 0.460 14.690 0.680 ;
        RECT 17.020 0.000 18.020 0.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 23.025 -4.020 23.455 -3.235 ;
      LAYER li1 ;
        RECT 20.180 -4.125 20.515 -3.385 ;
        RECT 23.095 -4.125 23.385 -3.400 ;
        RECT 20.090 -4.295 22.390 -4.125 ;
        RECT 23.010 -4.295 23.470 -4.125 ;
      LAYER met1 ;
        RECT 22.250 -3.970 23.220 -3.950 ;
        RECT 20.090 -4.450 23.470 -3.970 ;
        RECT 21.350 -5.250 22.350 -4.450 ;
    END
    PORT
      LAYER pwell ;
        RECT 28.095 -11.120 28.525 -10.335 ;
        RECT 15.605 -12.815 16.035 -12.030 ;
      LAYER li1 ;
        RECT 7.870 -11.235 8.100 -10.415 ;
        RECT 11.315 -11.235 11.625 -10.435 ;
        RECT 15.690 -11.235 15.920 -10.415 ;
        RECT 18.910 -11.235 19.140 -10.415 ;
        RECT 22.360 -11.235 22.615 -10.745 ;
        RECT 26.730 -11.235 26.960 -10.415 ;
        RECT 28.165 -11.225 28.455 -10.500 ;
        RECT 7.550 -11.405 8.930 -11.235 ;
        RECT 11.230 -11.405 12.610 -11.235 ;
        RECT 15.370 -11.405 16.750 -11.235 ;
        RECT 18.590 -11.405 19.970 -11.235 ;
        RECT 22.270 -11.405 24.110 -11.235 ;
        RECT 26.410 -11.405 27.790 -11.235 ;
        RECT 28.080 -11.395 28.540 -11.225 ;
        RECT 10.770 -11.795 12.150 -11.625 ;
        RECT 11.755 -12.595 12.065 -11.795 ;
        RECT 14.000 -11.855 15.380 -11.685 ;
        RECT 14.985 -12.655 15.295 -11.855 ;
        RECT 15.590 -11.925 16.050 -11.755 ;
        RECT 15.675 -12.650 15.965 -11.925 ;
      LAYER met1 ;
        RECT 27.900 -11.070 28.200 -11.050 ;
        RECT 27.900 -11.080 28.540 -11.070 ;
        RECT 7.550 -11.220 28.540 -11.080 ;
        RECT 7.360 -11.550 28.540 -11.220 ;
        RECT 7.360 -11.560 28.520 -11.550 ;
        RECT 7.360 -11.900 28.010 -11.560 ;
        RECT 10.770 -11.950 12.150 -11.900 ;
        RECT 14.000 -12.010 15.380 -11.900 ;
        RECT 15.590 -12.080 16.050 -11.900 ;
        RECT 25.000 -12.400 26.000 -11.900 ;
    END
  END VGND
  PIN f_vco
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 6.900 -10.005 8.170 -10.000 ;
        RECT 6.900 -10.200 8.200 -10.005 ;
        RECT 7.870 -10.245 8.200 -10.200 ;
      LAYER met1 ;
        RECT 3.250 -10.000 4.250 -9.700 ;
        RECT 4.820 -10.000 5.080 -9.940 ;
        RECT 3.250 -10.200 5.080 -10.000 ;
        RECT 3.250 -10.700 4.250 -10.200 ;
        RECT 4.820 -10.260 5.080 -10.200 ;
        RECT 6.190 -10.000 6.510 -9.970 ;
        RECT 6.870 -10.000 7.130 -9.940 ;
        RECT 6.190 -10.200 7.130 -10.000 ;
        RECT 6.190 -10.230 6.510 -10.200 ;
        RECT 6.870 -10.260 7.130 -10.200 ;
      LAYER met2 ;
        RECT 4.790 -10.000 5.110 -9.970 ;
        RECT 6.220 -10.000 6.480 -9.940 ;
        RECT 4.790 -10.200 6.480 -10.000 ;
        RECT 4.790 -10.230 5.110 -10.200 ;
        RECT 6.220 -10.260 6.480 -10.200 ;
    END
  END f_vco
  OBS
      LAYER pwell ;
        RECT 6.840 1.705 7.770 2.615 ;
        RECT 10.335 1.705 11.685 2.615 ;
        RECT 14.660 1.705 15.590 2.615 ;
        RECT 17.880 1.705 18.810 2.615 ;
        RECT 21.355 1.705 23.185 2.615 ;
        RECT 25.700 1.705 26.630 2.615 ;
        RECT 6.840 1.685 6.945 1.705 ;
        RECT 6.775 1.515 6.945 1.685 ;
        RECT 10.450 1.515 10.620 1.705 ;
        RECT 14.660 1.685 14.765 1.705 ;
        RECT 17.880 1.685 17.985 1.705 ;
        RECT 14.595 1.515 14.765 1.685 ;
        RECT 17.815 1.515 17.985 1.685 ;
        RECT 21.500 1.515 21.670 1.705 ;
        RECT 25.700 1.685 25.805 1.705 ;
        RECT 25.635 1.515 25.805 1.685 ;
        RECT 9.600 0.545 9.770 0.735 ;
        RECT 13.450 0.595 13.620 0.785 ;
        RECT 9.485 -0.365 10.835 0.545 ;
        RECT 13.335 -0.315 14.685 0.595 ;
        RECT 20.095 -4.105 22.385 -3.195 ;
        RECT 20.240 -4.295 20.410 -4.105 ;
        RECT 7.760 -11.215 8.690 -10.305 ;
        RECT 11.255 -11.215 12.605 -10.305 ;
        RECT 15.580 -11.215 16.510 -10.305 ;
        RECT 18.800 -11.215 19.730 -10.305 ;
        RECT 22.275 -11.215 24.105 -10.305 ;
        RECT 26.620 -11.215 27.550 -10.305 ;
        RECT 7.760 -11.235 7.865 -11.215 ;
        RECT 7.695 -11.405 7.865 -11.235 ;
        RECT 11.370 -11.405 11.540 -11.215 ;
        RECT 15.580 -11.235 15.685 -11.215 ;
        RECT 18.800 -11.235 18.905 -11.215 ;
        RECT 15.515 -11.405 15.685 -11.235 ;
        RECT 18.735 -11.405 18.905 -11.235 ;
        RECT 22.420 -11.405 22.590 -11.215 ;
        RECT 26.620 -11.235 26.725 -11.215 ;
        RECT 26.555 -11.405 26.725 -11.235 ;
        RECT 11.840 -11.815 12.010 -11.625 ;
        RECT 10.775 -12.725 12.125 -11.815 ;
        RECT 15.070 -11.875 15.240 -11.685 ;
        RECT 14.005 -12.785 15.355 -11.875 ;
      LAYER li1 ;
        RECT 7.350 3.085 7.680 4.065 ;
        RECT 10.845 3.085 11.175 4.065 ;
        RECT 13.175 3.475 13.925 3.730 ;
        RECT 7.450 2.900 7.680 3.085 ;
        RECT 10.405 2.900 10.740 2.925 ;
        RECT 7.450 2.700 10.740 2.900 ;
        RECT 7.450 2.485 7.680 2.700 ;
        RECT 10.405 2.655 10.740 2.700 ;
        RECT 7.350 1.855 7.680 2.485 ;
        RECT 10.910 2.485 11.080 3.085 ;
        RECT 11.250 2.900 11.585 2.925 ;
        RECT 13.700 2.900 13.890 3.475 ;
        RECT 15.170 3.085 15.500 4.065 ;
        RECT 18.390 3.085 18.720 4.065 ;
        RECT 14.770 2.900 15.100 2.915 ;
        RECT 11.250 2.700 12.350 2.900 ;
        RECT 13.700 2.700 15.100 2.900 ;
        RECT 11.250 2.675 11.585 2.700 ;
        RECT 10.910 2.200 11.605 2.485 ;
        RECT 13.700 2.200 13.900 2.700 ;
        RECT 14.770 2.675 15.100 2.700 ;
        RECT 15.270 2.900 15.500 3.085 ;
        RECT 17.990 2.900 18.320 2.915 ;
        RECT 15.270 2.700 18.320 2.900 ;
        RECT 15.270 2.485 15.500 2.700 ;
        RECT 17.990 2.675 18.320 2.700 ;
        RECT 18.490 2.850 18.720 3.085 ;
        RECT 19.900 2.850 20.100 3.800 ;
        RECT 21.865 3.265 22.195 4.065 ;
        RECT 22.765 3.265 23.095 4.065 ;
        RECT 21.865 3.095 23.095 3.265 ;
        RECT 24.400 3.250 25.050 3.450 ;
        RECT 21.460 2.850 21.680 2.925 ;
        RECT 18.490 2.650 20.100 2.850 ;
        RECT 20.750 2.650 21.680 2.850 ;
        RECT 18.490 2.485 18.720 2.650 ;
        RECT 10.910 2.000 13.900 2.200 ;
        RECT 10.910 1.855 11.605 2.000 ;
        RECT 15.170 1.855 15.500 2.485 ;
        RECT 18.390 1.855 18.720 2.485 ;
        RECT 20.750 1.800 20.950 2.650 ;
        RECT 21.460 2.345 21.680 2.650 ;
        RECT 21.865 2.195 22.045 3.095 ;
        RECT 22.215 2.365 22.590 2.925 ;
        RECT 22.795 2.900 23.105 2.925 ;
        RECT 24.850 2.900 25.050 3.250 ;
        RECT 26.210 3.085 26.540 4.065 ;
        RECT 25.810 2.900 26.140 2.915 ;
        RECT 22.795 2.650 24.100 2.900 ;
        RECT 24.850 2.700 26.140 2.900 ;
        RECT 22.795 2.595 23.105 2.650 ;
        RECT 22.765 2.195 23.095 2.425 ;
        RECT 23.855 2.405 24.050 2.650 ;
        RECT 21.865 2.150 23.095 2.195 ;
        RECT 24.850 2.150 25.050 2.700 ;
        RECT 25.810 2.675 26.140 2.700 ;
        RECT 26.310 2.900 26.540 3.085 ;
        RECT 26.310 2.700 27.950 2.900 ;
        RECT 26.310 2.485 26.540 2.700 ;
        RECT 21.865 1.950 25.050 2.150 ;
        RECT 21.865 1.855 23.095 1.950 ;
        RECT 26.210 1.855 26.540 2.485 ;
        RECT 10.060 0.250 10.755 0.395 ;
        RECT 10.060 0.050 11.750 0.250 ;
        RECT 13.910 0.200 14.605 0.445 ;
        RECT 10.060 -0.235 10.755 0.050 ;
        RECT 13.910 0.000 15.900 0.200 ;
        RECT 13.910 -0.185 14.605 0.000 ;
        RECT 9.555 -0.450 9.890 -0.405 ;
        RECT 8.400 -0.650 9.890 -0.450 ;
        RECT 9.555 -0.675 9.890 -0.650 ;
        RECT 10.060 -0.835 10.230 -0.235 ;
        RECT 13.405 -0.400 13.740 -0.355 ;
        RECT 10.400 -0.450 10.735 -0.425 ;
        RECT 10.400 -0.650 12.350 -0.450 ;
        RECT 12.650 -0.600 13.740 -0.400 ;
        RECT 13.405 -0.625 13.740 -0.600 ;
        RECT 10.400 -0.675 10.735 -0.650 ;
        RECT 9.995 -1.815 10.325 -0.835 ;
        RECT 11.425 -0.950 11.625 -0.650 ;
        RECT 13.910 -0.785 14.080 -0.185 ;
        RECT 14.250 -0.415 14.585 -0.375 ;
        RECT 14.250 -0.585 15.185 -0.415 ;
        RECT 14.250 -0.625 14.585 -0.585 ;
        RECT 13.845 -1.765 14.175 -0.785 ;
        RECT 18.600 -2.250 18.800 -1.600 ;
        RECT 18.600 -2.450 19.550 -2.250 ;
        RECT 20.605 -2.545 20.935 -1.745 ;
        RECT 21.475 -2.545 21.805 -1.745 ;
        RECT 20.605 -2.715 21.885 -2.545 ;
        RECT 17.640 -2.950 19.760 -2.940 ;
        RECT 20.200 -2.950 20.485 -2.885 ;
        RECT 17.640 -3.150 20.500 -2.950 ;
        RECT 17.640 -3.160 19.760 -3.150 ;
        RECT 20.200 -3.215 20.485 -3.150 ;
        RECT 20.685 -3.215 21.065 -2.885 ;
        RECT 21.235 -3.215 21.545 -2.885 ;
        RECT 18.700 -3.800 19.800 -3.600 ;
        RECT 18.705 -5.145 18.895 -3.800 ;
        RECT 20.685 -3.910 20.900 -3.215 ;
        RECT 21.235 -3.385 21.440 -3.215 ;
        RECT 21.715 -3.385 21.885 -2.715 ;
        RECT 22.065 -2.950 22.305 -2.545 ;
        RECT 22.065 -3.150 24.850 -2.950 ;
        RECT 22.065 -3.215 22.305 -3.150 ;
        RECT 21.090 -3.910 21.440 -3.385 ;
        RECT 21.610 -3.955 22.305 -3.385 ;
        RECT 8.270 -9.835 8.600 -8.855 ;
        RECT 11.765 -9.835 12.095 -8.855 ;
        RECT 16.090 -9.835 16.420 -8.855 ;
        RECT 19.310 -9.835 19.640 -8.855 ;
        RECT 8.370 -10.050 8.600 -9.835 ;
        RECT 11.325 -10.050 11.660 -9.995 ;
        RECT 8.370 -10.250 11.660 -10.050 ;
        RECT 8.370 -10.435 8.600 -10.250 ;
        RECT 11.325 -10.265 11.660 -10.250 ;
        RECT 8.270 -11.065 8.600 -10.435 ;
        RECT 11.830 -10.435 12.000 -9.835 ;
        RECT 12.170 -10.000 12.505 -9.995 ;
        RECT 16.190 -10.000 16.420 -9.835 ;
        RECT 12.170 -10.200 13.250 -10.000 ;
        RECT 14.850 -10.005 15.950 -10.000 ;
        RECT 16.190 -10.005 19.150 -10.000 ;
        RECT 14.850 -10.200 16.020 -10.005 ;
        RECT 12.170 -10.245 12.505 -10.200 ;
        RECT 11.830 -10.700 12.525 -10.435 ;
        RECT 14.200 -10.700 14.400 -10.250 ;
        RECT 14.850 -10.700 15.050 -10.200 ;
        RECT 15.690 -10.245 16.020 -10.200 ;
        RECT 16.190 -10.200 19.240 -10.005 ;
        RECT 16.190 -10.435 16.420 -10.200 ;
        RECT 18.910 -10.245 19.240 -10.200 ;
        RECT 19.410 -10.050 19.640 -9.835 ;
        RECT 22.785 -9.655 23.115 -8.855 ;
        RECT 23.685 -9.655 24.015 -8.855 ;
        RECT 22.785 -9.825 24.015 -9.655 ;
        RECT 22.380 -10.050 22.600 -9.995 ;
        RECT 19.410 -10.250 21.500 -10.050 ;
        RECT 21.700 -10.250 22.600 -10.050 ;
        RECT 19.410 -10.435 19.640 -10.250 ;
        RECT 11.830 -10.900 15.050 -10.700 ;
        RECT 11.830 -11.065 12.525 -10.900 ;
        RECT 16.090 -11.065 16.420 -10.435 ;
        RECT 19.310 -11.065 19.640 -10.435 ;
        RECT 22.380 -10.575 22.600 -10.250 ;
        RECT 22.785 -10.725 22.965 -9.825 ;
        RECT 27.130 -9.835 27.460 -8.855 ;
        RECT 23.135 -10.555 23.510 -9.995 ;
        RECT 23.715 -10.065 24.025 -9.995 ;
        RECT 25.500 -10.065 26.350 -10.050 ;
        RECT 26.730 -10.065 27.060 -10.005 ;
        RECT 23.715 -10.235 24.780 -10.065 ;
        RECT 25.500 -10.235 27.060 -10.065 ;
        RECT 23.715 -10.325 24.025 -10.235 ;
        RECT 25.500 -10.250 26.350 -10.235 ;
        RECT 26.730 -10.245 27.060 -10.235 ;
        RECT 27.230 -10.050 27.460 -9.835 ;
        RECT 23.685 -10.725 24.015 -10.495 ;
        RECT 22.785 -10.750 24.015 -10.725 ;
        RECT 26.150 -10.750 26.350 -10.250 ;
        RECT 27.230 -10.250 29.900 -10.050 ;
        RECT 27.230 -10.435 27.460 -10.250 ;
        RECT 22.785 -10.950 26.350 -10.750 ;
        RECT 22.785 -11.065 24.015 -10.950 ;
        RECT 27.130 -11.065 27.460 -10.435 ;
        RECT 10.855 -12.350 11.550 -11.965 ;
        RECT 14.085 -12.200 14.780 -12.025 ;
        RECT 9.800 -12.550 11.550 -12.350 ;
        RECT 10.855 -12.595 11.550 -12.550 ;
        RECT 10.875 -12.865 11.210 -12.785 ;
        RECT 9.565 -13.035 11.210 -12.865 ;
        RECT 11.380 -13.195 11.550 -12.595 ;
        RECT 12.350 -12.400 14.780 -12.200 ;
        RECT 11.720 -12.800 12.055 -12.765 ;
        RECT 12.350 -12.800 12.550 -12.400 ;
        RECT 11.720 -13.000 12.550 -12.800 ;
        RECT 11.720 -13.035 12.055 -13.000 ;
        RECT 11.285 -14.175 11.615 -13.195 ;
        RECT 12.900 -13.700 13.100 -12.400 ;
        RECT 14.085 -12.655 14.780 -12.400 ;
        RECT 14.105 -12.865 14.440 -12.845 ;
        RECT 13.565 -13.035 14.440 -12.865 ;
        RECT 14.105 -13.095 14.440 -13.035 ;
        RECT 14.610 -13.255 14.780 -12.655 ;
        RECT 14.950 -12.850 15.285 -12.825 ;
        RECT 14.950 -13.050 16.700 -12.850 ;
        RECT 14.950 -13.095 15.285 -13.050 ;
        RECT 14.515 -14.235 14.845 -13.255 ;
      LAYER met1 ;
        RECT 12.120 6.550 12.380 6.610 ;
        RECT 24.340 6.550 24.660 6.580 ;
        RECT 12.120 6.350 24.660 6.550 ;
        RECT 12.120 6.290 12.380 6.350 ;
        RECT 24.340 6.320 24.660 6.350 ;
        RECT 33.450 5.670 33.770 5.700 ;
        RECT 32.800 5.470 33.770 5.670 ;
        RECT 12.090 3.620 12.410 3.880 ;
        RECT 24.370 3.840 24.630 4.160 ;
        RECT 19.840 3.800 20.160 3.830 ;
        RECT 12.150 2.915 12.350 3.620 ;
        RECT 13.150 3.100 13.450 3.780 ;
        RECT 19.840 3.600 22.450 3.800 ;
        RECT 19.840 3.570 20.160 3.600 ;
        RECT 12.105 2.685 12.395 2.915 ;
        RECT 13.120 2.800 13.480 3.100 ;
        RECT 22.250 2.845 22.450 3.600 ;
        RECT 24.400 3.510 24.600 3.840 ;
        RECT 24.370 3.190 24.630 3.510 ;
        RECT 27.670 2.900 27.930 2.960 ;
        RECT 32.800 2.900 33.000 5.470 ;
        RECT 33.450 5.440 33.770 5.470 ;
        RECT 34.730 5.670 34.990 5.730 ;
        RECT 34.730 5.470 35.860 5.670 ;
        RECT 34.730 5.410 34.990 5.470 ;
        RECT 22.235 2.555 22.465 2.845 ;
        RECT 27.670 2.700 33.000 2.900 ;
        RECT 23.825 2.630 24.085 2.665 ;
        RECT 27.670 2.640 27.930 2.700 ;
        RECT 23.795 2.375 24.110 2.630 ;
        RECT 23.825 2.345 24.085 2.375 ;
        RECT 19.640 2.000 19.960 2.030 ;
        RECT 20.705 2.000 20.995 2.015 ;
        RECT 19.640 1.800 20.995 2.000 ;
        RECT 19.640 1.770 19.960 1.800 ;
        RECT 20.705 1.785 20.995 1.800 ;
        RECT 11.520 -0.010 11.780 0.310 ;
        RECT 12.120 -0.010 12.380 0.310 ;
        RECT 14.940 0.170 15.260 0.430 ;
        RECT 12.150 -0.390 12.350 -0.010 ;
        RECT 8.355 -0.665 8.645 -0.435 ;
        RECT 8.400 -3.550 8.600 -0.665 ;
        RECT 11.410 -0.720 11.670 -0.690 ;
        RECT 12.120 -0.710 12.380 -0.390 ;
        RECT 12.620 -0.660 12.880 -0.340 ;
        RECT 15.020 -0.355 15.180 0.170 ;
        RECT 15.670 -0.060 15.930 0.260 ;
        RECT 19.640 0.170 19.960 0.430 ;
        RECT 14.985 -0.645 15.215 -0.355 ;
        RECT 11.380 -0.980 11.670 -0.720 ;
        RECT 11.410 -1.010 11.670 -0.980 ;
        RECT 11.445 -1.655 11.765 -1.615 ;
        RECT 12.660 -1.655 12.845 -0.660 ;
        RECT 11.445 -1.840 12.845 -1.655 ;
        RECT 11.445 -1.875 11.765 -1.840 ;
        RECT 15.700 -3.550 15.900 -0.060 ;
        RECT 19.700 -0.150 19.900 0.170 ;
        RECT 19.700 -0.350 24.850 -0.150 ;
        RECT 18.570 -1.010 18.830 -0.690 ;
        RECT 18.600 -1.555 18.800 -1.010 ;
        RECT 18.585 -1.845 18.815 -1.555 ;
        RECT 19.320 -2.250 19.580 -2.190 ;
        RECT 19.320 -2.450 20.950 -2.250 ;
        RECT 19.320 -2.510 19.580 -2.450 ;
        RECT 20.750 -2.905 20.950 -2.450 ;
        RECT 24.650 -2.905 24.850 -0.350 ;
        RECT 17.605 -3.165 17.895 -2.935 ;
        RECT 8.400 -3.750 15.900 -3.550 ;
        RECT 11.450 -4.275 11.770 -4.015 ;
        RECT 11.520 -5.545 11.705 -4.275 ;
        RECT 13.640 -4.790 13.960 -4.770 ;
        RECT 17.640 -4.790 17.860 -3.165 ;
        RECT 20.735 -3.195 20.965 -2.905 ;
        RECT 24.635 -3.195 24.865 -2.905 ;
        RECT 21.710 -3.500 22.000 -3.475 ;
        RECT 22.425 -3.500 22.685 -3.435 ;
        RECT 19.570 -3.600 19.830 -3.540 ;
        RECT 21.105 -3.600 21.395 -3.585 ;
        RECT 19.570 -3.800 21.395 -3.600 ;
        RECT 21.710 -3.685 22.685 -3.500 ;
        RECT 21.710 -3.705 22.000 -3.685 ;
        RECT 22.425 -3.755 22.685 -3.685 ;
        RECT 19.570 -3.860 19.830 -3.800 ;
        RECT 21.105 -3.815 21.395 -3.800 ;
        RECT 13.640 -5.010 17.860 -4.790 ;
        RECT 18.655 -4.955 18.945 -4.935 ;
        RECT 20.640 -4.955 20.960 -4.920 ;
        RECT 13.640 -5.030 13.960 -5.010 ;
        RECT 18.655 -5.145 20.960 -4.955 ;
        RECT 18.655 -5.165 18.945 -5.145 ;
        RECT 20.640 -5.180 20.960 -5.145 ;
        RECT 23.140 -5.545 23.460 -5.505 ;
        RECT 11.520 -5.730 23.460 -5.545 ;
        RECT 11.520 -7.405 11.705 -5.730 ;
        RECT 23.140 -5.765 23.460 -5.730 ;
        RECT 5.660 -7.590 11.705 -7.405 ;
        RECT 13.050 -6.600 25.700 -6.400 ;
        RECT 13.050 -7.490 13.250 -6.600 ;
        RECT 25.500 -7.470 25.700 -6.600 ;
        RECT 5.665 -14.570 5.835 -7.590 ;
        RECT 13.020 -7.810 13.280 -7.490 ;
        RECT 25.440 -7.730 25.760 -7.470 ;
        RECT 12.990 -9.330 13.310 -9.070 ;
        RECT 21.250 -9.250 23.450 -9.050 ;
        RECT 13.050 -9.985 13.250 -9.330 ;
        RECT 14.170 -9.580 14.430 -9.260 ;
        RECT 13.640 -9.800 13.960 -9.770 ;
        RECT 14.200 -9.800 14.400 -9.580 ;
        RECT 13.005 -10.215 13.295 -9.985 ;
        RECT 13.640 -10.000 14.400 -9.800 ;
        RECT 13.640 -10.030 13.960 -10.000 ;
        RECT 14.200 -10.235 14.400 -10.000 ;
        RECT 21.250 -10.020 21.450 -9.250 ;
        RECT 14.155 -10.465 14.445 -10.235 ;
        RECT 21.190 -10.280 21.510 -10.020 ;
        RECT 21.655 -10.265 21.945 -10.035 ;
        RECT 23.250 -10.055 23.450 -9.250 ;
        RECT 24.535 -9.330 24.855 -9.070 ;
        RECT 25.470 -9.310 25.730 -8.990 ;
        RECT 24.610 -10.005 24.780 -9.330 ;
        RECT 25.500 -9.990 25.700 -9.310 ;
        RECT 21.700 -10.620 21.900 -10.265 ;
        RECT 23.235 -10.345 23.465 -10.055 ;
        RECT 24.580 -10.295 24.810 -10.005 ;
        RECT 25.470 -10.310 25.730 -9.990 ;
        RECT 29.670 -10.050 29.930 -9.990 ;
        RECT 35.170 -10.050 35.490 -10.020 ;
        RECT 29.670 -10.250 35.490 -10.050 ;
        RECT 29.670 -10.310 29.930 -10.250 ;
        RECT 35.170 -10.280 35.490 -10.250 ;
        RECT 36.530 -10.050 36.790 -9.990 ;
        RECT 37.050 -10.050 37.250 -8.160 ;
        RECT 36.530 -10.250 37.250 -10.050 ;
        RECT 36.530 -10.310 36.790 -10.250 ;
        RECT 21.640 -10.880 21.960 -10.620 ;
        RECT 9.770 -12.610 10.030 -12.290 ;
        RECT 13.490 -12.480 13.810 -12.220 ;
        RECT 16.470 -12.410 16.730 -12.090 ;
        RECT 13.565 -12.805 13.735 -12.480 ;
        RECT 9.505 -13.065 9.795 -12.835 ;
        RECT 9.570 -14.570 9.730 -13.065 ;
        RECT 13.535 -13.095 13.765 -12.805 ;
        RECT 16.500 -12.820 16.700 -12.410 ;
        RECT 20.670 -12.460 20.930 -12.140 ;
        RECT 16.440 -13.080 16.760 -12.820 ;
        RECT 12.840 -13.500 13.160 -13.470 ;
        RECT 20.700 -13.500 20.900 -12.460 ;
        RECT 21.670 -12.560 21.930 -12.240 ;
        RECT 21.700 -13.500 21.900 -12.560 ;
        RECT 12.840 -13.700 21.900 -13.500 ;
        RECT 12.840 -13.730 13.160 -13.700 ;
        RECT 5.665 -14.730 9.730 -14.570 ;
        RECT 5.665 -14.735 5.835 -14.730 ;
      LAYER met2 ;
        RECT 12.090 6.320 12.410 6.580 ;
        RECT 12.150 3.910 12.350 6.320 ;
        RECT 24.370 6.290 24.630 6.610 ;
        RECT 24.400 4.130 24.600 6.290 ;
        RECT 33.480 5.670 33.740 5.730 ;
        RECT 34.700 5.670 35.020 5.700 ;
        RECT 33.480 5.470 35.020 5.670 ;
        RECT 33.480 5.410 33.740 5.470 ;
        RECT 34.700 5.440 35.020 5.470 ;
        RECT 12.120 3.590 12.380 3.910 ;
        RECT 24.340 3.870 24.660 4.130 ;
        RECT 12.110 1.850 12.390 1.885 ;
        RECT 13.150 1.850 13.450 3.130 ;
        RECT 23.795 2.375 24.115 2.635 ;
        RECT 12.100 1.550 13.450 1.850 ;
        RECT 19.670 1.740 19.930 2.060 ;
        RECT 12.110 1.515 12.390 1.550 ;
        RECT 19.700 1.200 19.900 1.740 ;
        RECT 11.550 1.000 19.900 1.200 ;
        RECT 11.550 0.280 11.750 1.000 ;
        RECT 15.000 0.460 15.200 1.000 ;
        RECT 19.700 0.460 19.900 1.000 ;
        RECT 12.100 0.280 12.400 0.345 ;
        RECT 11.490 0.020 11.810 0.280 ;
        RECT 12.090 0.020 12.410 0.280 ;
        RECT 14.970 0.140 15.230 0.460 ;
        RECT 19.670 0.140 19.930 0.460 ;
        RECT 12.100 -0.045 12.400 0.020 ;
        RECT 23.860 -0.495 24.055 2.375 ;
        RECT 11.380 -0.750 11.700 -0.720 ;
        RECT 18.540 -0.750 18.860 -0.720 ;
        RECT 11.380 -0.950 18.860 -0.750 ;
        RECT 11.380 -0.980 11.700 -0.950 ;
        RECT 18.540 -0.980 18.860 -0.950 ;
        RECT 11.475 -1.905 11.735 -1.585 ;
        RECT 11.515 -3.985 11.700 -1.905 ;
        RECT 22.395 -3.505 22.715 -3.465 ;
        RECT 23.865 -3.505 24.050 -0.495 ;
        RECT 22.395 -3.690 24.050 -3.505 ;
        RECT 22.395 -3.725 22.715 -3.690 ;
        RECT 11.480 -4.305 11.740 -3.985 ;
        RECT 13.670 -5.060 13.930 -4.740 ;
        RECT 13.690 -7.360 13.910 -5.060 ;
        RECT 20.670 -5.210 20.930 -4.890 ;
        RECT 12.990 -7.780 13.310 -7.520 ;
        RECT 13.050 -9.040 13.250 -7.780 ;
        RECT 13.020 -9.360 13.280 -9.040 ;
        RECT 13.700 -9.740 13.900 -7.360 ;
        RECT 14.140 -9.320 14.460 -9.290 ;
        RECT 14.760 -9.320 16.700 -9.300 ;
        RECT 14.140 -9.500 16.700 -9.320 ;
        RECT 14.140 -9.520 14.910 -9.500 ;
        RECT 14.140 -9.550 14.460 -9.520 ;
        RECT 13.670 -10.060 13.930 -9.740 ;
        RECT 9.800 -11.500 13.750 -11.300 ;
        RECT 9.800 -12.320 10.000 -11.500 ;
        RECT 13.550 -12.190 13.750 -11.500 ;
        RECT 16.500 -12.120 16.700 -9.500 ;
        RECT 9.740 -12.580 10.060 -12.320 ;
        RECT 13.520 -12.510 13.780 -12.190 ;
        RECT 16.440 -12.380 16.760 -12.120 ;
        RECT 20.700 -12.170 20.900 -5.210 ;
        RECT 23.170 -5.540 23.430 -5.475 ;
        RECT 23.865 -5.540 24.050 -3.690 ;
        RECT 23.170 -5.725 24.050 -5.540 ;
        RECT 23.170 -5.795 23.430 -5.725 ;
        RECT 23.865 -7.305 24.050 -5.725 ;
        RECT 23.865 -7.490 24.790 -7.305 ;
        RECT 24.610 -9.040 24.780 -7.490 ;
        RECT 25.470 -7.760 25.730 -7.440 ;
        RECT 25.500 -9.020 25.700 -7.760 ;
        RECT 24.565 -9.360 24.825 -9.040 ;
        RECT 25.440 -9.280 25.760 -9.020 ;
        RECT 35.200 -10.050 35.460 -9.990 ;
        RECT 36.500 -10.050 36.820 -10.020 ;
        RECT 35.200 -10.250 36.820 -10.050 ;
        RECT 35.200 -10.310 35.460 -10.250 ;
        RECT 36.500 -10.280 36.820 -10.250 ;
        RECT 21.670 -10.910 21.930 -10.590 ;
        RECT 20.640 -12.430 20.960 -12.170 ;
        RECT 21.700 -12.270 21.900 -10.910 ;
        RECT 21.640 -12.530 21.960 -12.270 ;
      LAYER met3 ;
        RECT 12.085 1.535 12.415 1.865 ;
        RECT 12.100 0.325 12.400 1.535 ;
        RECT 12.075 -0.025 12.425 0.325 ;
  END
END pfd_lay
MACRO cp
  CLASS BLOCK ;
  FOREIGN cp ;
  ORIGIN 327.630 5.220 ;
  SIZE 586.465 BY 447.730 ;
  PIN up
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.185 27.370 2.515 27.540 ;
        RECT 2.185 26.190 2.515 26.360 ;
        RECT 2.205 24.430 2.535 24.600 ;
        RECT 2.205 23.460 2.535 23.630 ;
        RECT 18.445 19.800 18.775 19.970 ;
        RECT 18.445 18.620 18.775 18.790 ;
      LAYER met1 ;
        RECT -0.380 27.350 2.530 27.580 ;
        RECT -0.380 26.375 -0.150 27.350 ;
        RECT 2.205 27.340 2.495 27.350 ;
        RECT 2.205 26.375 2.495 26.390 ;
        RECT -0.380 26.160 2.495 26.375 ;
        RECT -0.380 26.145 2.485 26.160 ;
        RECT -2.430 25.490 -1.430 25.860 ;
        RECT -0.380 25.490 -0.150 26.145 ;
        RECT -2.430 25.270 -0.150 25.490 ;
        RECT -2.430 24.860 -1.430 25.270 ;
        RECT -0.940 18.200 -0.720 25.270 ;
        RECT -0.380 24.665 -0.150 25.270 ;
        RECT -0.380 24.435 2.525 24.665 ;
        RECT -0.380 23.645 -0.150 24.435 ;
        RECT 2.225 24.400 2.515 24.435 ;
        RECT 2.225 23.645 2.515 23.660 ;
        RECT -0.380 23.415 2.525 23.645 ;
        RECT 16.020 20.000 18.740 20.010 ;
        RECT 16.020 19.790 18.755 20.000 ;
        RECT 16.020 18.770 16.240 19.790 ;
        RECT 18.465 19.770 18.755 19.790 ;
        RECT 18.465 18.770 18.755 18.820 ;
        RECT 16.000 18.550 18.780 18.770 ;
        RECT 1.540 18.200 1.860 18.220 ;
        RECT -0.940 17.980 1.860 18.200 ;
        RECT 1.540 17.960 1.860 17.980 ;
        RECT 3.070 18.200 3.330 18.250 ;
        RECT 5.880 18.200 6.200 18.220 ;
        RECT 3.070 17.980 6.200 18.200 ;
        RECT 3.070 17.930 3.330 17.980 ;
        RECT 5.880 17.960 6.200 17.980 ;
        RECT 7.730 18.200 7.990 18.250 ;
        RECT 16.000 18.200 16.220 18.550 ;
        RECT 7.730 17.980 16.220 18.200 ;
        RECT 7.730 17.930 7.990 17.980 ;
      LAYER met2 ;
        RECT 1.570 18.200 1.830 18.250 ;
        RECT 3.040 18.200 3.360 18.220 ;
        RECT 1.570 17.980 3.360 18.200 ;
        RECT 1.570 17.930 1.830 17.980 ;
        RECT 3.040 17.960 3.360 17.980 ;
        RECT 5.910 18.200 6.170 18.250 ;
        RECT 7.700 18.200 8.020 18.220 ;
        RECT 5.910 17.980 8.020 18.200 ;
        RECT 5.910 17.930 6.170 17.980 ;
        RECT 7.700 17.960 8.020 17.980 ;
    END
  END up
  PIN vctrl
    ANTENNADIFFAREA 0.278400 ;
    PORT
      LAYER li1 ;
        RECT 57.600 37.150 57.920 38.965 ;
        RECT 57.520 36.980 58.000 37.150 ;
        RECT 26.650 26.495 26.820 27.075 ;
        RECT 33.920 12.680 34.090 13.140 ;
      LAYER met1 ;
        RECT 74.680 98.020 85.450 98.460 ;
        RECT 57.570 36.920 57.950 39.025 ;
        RECT 57.600 35.870 57.920 36.920 ;
        RECT 57.600 35.520 57.900 35.870 ;
        RECT 57.560 35.080 57.900 35.520 ;
        RECT 57.600 34.680 57.900 35.080 ;
        RECT 57.600 29.720 57.920 34.680 ;
        RECT 36.710 29.400 57.920 29.720 ;
        RECT 26.620 26.920 26.850 27.055 ;
        RECT 26.620 26.710 28.210 26.920 ;
        RECT 26.620 26.515 26.850 26.710 ;
        RECT 28.000 21.020 28.210 26.710 ;
        RECT 36.710 21.020 37.030 29.400 ;
        RECT 74.680 24.120 75.120 98.020 ;
        RECT 40.530 23.680 75.120 24.120 ;
        RECT 40.530 21.020 40.970 23.680 ;
        RECT 44.960 21.020 45.960 21.230 ;
        RECT 27.970 20.660 45.960 21.020 ;
        RECT 28.000 14.295 28.210 20.660 ;
        RECT 44.960 20.210 45.960 20.660 ;
        RECT 32.790 14.295 33.110 14.320 ;
        RECT 28.000 14.085 33.110 14.295 ;
        RECT 32.790 14.060 33.110 14.085 ;
        RECT 32.790 13.005 33.110 13.030 ;
        RECT 33.890 13.005 34.120 13.120 ;
        RECT 32.790 12.795 34.120 13.005 ;
        RECT 32.790 12.770 33.110 12.795 ;
        RECT 33.890 12.700 34.120 12.795 ;
      LAYER met2 ;
        RECT 84.980 98.460 85.420 98.490 ;
        RECT 84.980 98.020 87.095 98.460 ;
        RECT 84.980 97.990 85.420 98.020 ;
        RECT 32.820 14.030 33.080 14.350 ;
        RECT 32.845 13.060 33.055 14.030 ;
        RECT 32.820 12.740 33.080 13.060 ;
      LAYER met3 ;
        RECT 255.990 183.000 256.570 183.520 ;
        RECT 256.020 179.195 256.540 183.000 ;
        RECT 255.995 178.685 256.565 179.195 ;
        RECT 256.020 178.680 256.540 178.685 ;
        RECT 86.585 98.460 87.075 98.485 ;
        RECT 86.585 98.020 88.890 98.460 ;
        RECT 86.585 97.995 87.075 98.020 ;
      LAYER met4 ;
        RECT 98.225 230.720 127.835 245.265 ;
        RECT 129.825 230.720 159.435 245.265 ;
        RECT 161.425 230.720 191.035 245.265 ;
        RECT 193.025 230.720 222.635 245.265 ;
        RECT 224.625 230.720 254.235 245.265 ;
        RECT 97.230 230.710 255.230 230.720 ;
        RECT 95.100 230.200 255.230 230.710 ;
        RECT 95.100 230.190 127.835 230.200 ;
        RECT 95.100 197.660 95.620 230.190 ;
        RECT 98.225 215.655 127.835 230.190 ;
        RECT 129.825 215.655 159.435 230.200 ;
        RECT 161.425 215.655 191.035 230.200 ;
        RECT 193.025 215.655 222.635 230.200 ;
        RECT 224.625 215.655 254.235 230.200 ;
        RECT 98.225 197.660 127.835 212.205 ;
        RECT 129.825 197.660 159.435 212.205 ;
        RECT 161.425 197.660 191.035 212.205 ;
        RECT 193.025 197.660 222.635 212.205 ;
        RECT 224.625 197.660 254.235 212.205 ;
        RECT 254.820 197.660 256.540 197.680 ;
        RECT 95.100 197.160 256.540 197.660 ;
        RECT 95.100 197.140 255.230 197.160 ;
        RECT 98.225 182.595 127.835 197.140 ;
        RECT 129.825 182.595 159.435 197.140 ;
        RECT 161.425 182.595 191.035 197.140 ;
        RECT 193.025 182.595 222.635 197.140 ;
        RECT 224.625 182.595 254.235 197.140 ;
        RECT 256.020 183.525 256.540 197.160 ;
        RECT 256.015 182.995 256.545 183.525 ;
        RECT 98.225 164.600 127.835 179.145 ;
        RECT 129.825 164.600 159.435 179.145 ;
        RECT 161.425 164.600 191.035 179.145 ;
        RECT 193.025 164.600 222.635 179.145 ;
        RECT 224.625 164.600 254.235 179.145 ;
        RECT 256.020 164.600 256.540 179.200 ;
        RECT 97.230 164.590 256.540 164.600 ;
        RECT 93.500 164.080 256.540 164.590 ;
        RECT 93.500 164.070 97.770 164.080 ;
        RECT 93.500 131.540 94.020 164.070 ;
        RECT 98.225 149.535 127.835 164.080 ;
        RECT 129.825 149.535 159.435 164.080 ;
        RECT 161.425 149.535 191.035 164.080 ;
        RECT 193.025 149.535 222.635 164.080 ;
        RECT 224.625 149.535 254.235 164.080 ;
        RECT 98.225 131.540 127.835 146.085 ;
        RECT 129.825 131.540 159.435 146.085 ;
        RECT 161.425 131.540 191.035 146.085 ;
        RECT 193.025 131.540 222.635 146.085 ;
        RECT 224.625 131.540 254.235 146.085 ;
        RECT 255.040 131.540 257.080 131.600 ;
        RECT 93.500 131.080 257.080 131.540 ;
        RECT 93.500 131.020 255.230 131.080 ;
        RECT 98.225 116.475 127.835 131.020 ;
        RECT 129.825 116.475 159.435 131.020 ;
        RECT 161.425 116.475 191.035 131.020 ;
        RECT 193.025 116.475 222.635 131.020 ;
        RECT 224.625 116.475 254.235 131.020 ;
        RECT 98.225 98.480 127.835 113.025 ;
        RECT 129.825 98.480 159.435 113.025 ;
        RECT 161.425 98.480 191.035 113.025 ;
        RECT 193.025 98.480 222.635 113.025 ;
        RECT 224.625 98.480 254.235 113.025 ;
        RECT 256.560 98.480 257.080 131.080 ;
        RECT 88.415 98.460 88.865 98.465 ;
        RECT 97.230 98.460 257.080 98.480 ;
        RECT 88.415 98.020 257.080 98.460 ;
        RECT 88.415 98.015 88.865 98.020 ;
        RECT 97.230 97.960 257.080 98.020 ;
        RECT 98.225 83.415 127.835 97.960 ;
        RECT 129.825 83.415 159.435 97.960 ;
        RECT 161.425 83.415 191.035 97.960 ;
        RECT 193.025 83.415 222.635 97.960 ;
        RECT 224.625 83.415 254.235 97.960 ;
    END
  END vctrl
  PIN VDD
    ANTENNAGATEAREA 0.345600 ;
    ANTENNADIFFAREA 33.939598 ;
    PORT
      LAYER nwell ;
        RECT -5.790 32.030 41.400 34.170 ;
        RECT 1.280 25.500 3.420 28.230 ;
        RECT 19.720 25.300 21.860 28.030 ;
        RECT 1.940 11.700 4.080 14.430 ;
      LAYER li1 ;
        RECT -5.610 33.820 41.220 33.990 ;
        RECT -5.610 32.380 -5.440 33.820 ;
        RECT -4.715 33.250 40.325 33.420 ;
        RECT 41.050 32.380 41.220 33.820 ;
        RECT -5.610 32.210 41.220 32.380 ;
        RECT 1.460 27.880 3.240 28.050 ;
        RECT 1.460 25.850 1.630 27.880 ;
        RECT 2.030 26.575 2.200 27.155 ;
        RECT 3.070 25.850 3.240 27.880 ;
        RECT 19.900 27.680 21.680 27.850 ;
        RECT 10.315 27.420 10.645 27.590 ;
        RECT 10.315 26.240 10.645 26.410 ;
        RECT 1.460 25.680 3.240 25.850 ;
        RECT 19.900 25.650 20.070 27.680 ;
        RECT 20.940 26.375 21.110 26.955 ;
        RECT 21.510 25.650 21.680 27.680 ;
        RECT 19.900 25.480 21.680 25.650 ;
        RECT 2.120 14.080 3.900 14.250 ;
        RECT 23.675 14.090 24.005 14.260 ;
        RECT 2.120 12.050 2.290 14.080 ;
        RECT 2.690 12.775 2.860 13.355 ;
        RECT 3.730 12.050 3.900 14.080 ;
        RECT 11.205 13.640 11.535 13.810 ;
        RECT 23.990 13.460 24.160 13.920 ;
        RECT 34.075 13.310 34.405 13.480 ;
        RECT 23.675 13.120 24.005 13.290 ;
        RECT 11.205 12.460 11.535 12.630 ;
        RECT 34.075 12.340 34.405 12.510 ;
        RECT 2.120 11.880 3.900 12.050 ;
      LAYER met1 ;
        RECT 39.120 34.745 39.350 34.790 ;
        RECT 39.120 34.515 41.795 34.745 ;
        RECT 39.120 33.450 39.350 34.515 ;
        RECT 41.565 34.050 41.795 34.515 ;
        RECT 22.150 33.220 40.220 33.450 ;
        RECT 40.980 32.230 41.990 34.050 ;
        RECT 41.425 30.905 41.755 32.230 ;
        RECT 33.755 30.575 41.755 30.905 ;
        RECT 19.220 30.195 19.550 30.210 ;
        RECT 26.535 30.195 26.865 30.225 ;
        RECT 33.755 30.195 34.085 30.575 ;
        RECT 8.850 29.720 9.850 30.110 ;
        RECT -3.750 29.370 9.850 29.720 ;
        RECT -3.750 15.365 -3.400 29.370 ;
        RECT 8.850 29.000 9.850 29.370 ;
        RECT 19.220 29.865 22.815 30.195 ;
        RECT 26.535 29.865 34.085 30.195 ;
        RECT 19.220 29.260 19.550 29.865 ;
        RECT 26.535 29.835 26.865 29.865 ;
        RECT 19.050 29.000 19.550 29.260 ;
        RECT 1.400 28.970 19.550 29.000 ;
        RECT 1.400 28.450 19.630 28.970 ;
        RECT 0.640 28.070 0.960 28.100 ;
        RECT 1.490 28.070 3.350 28.450 ;
        RECT 0.640 27.880 3.350 28.070 ;
        RECT 0.640 27.870 3.130 27.880 ;
        RECT 0.640 27.840 0.960 27.870 ;
        RECT 1.570 27.850 3.130 27.870 ;
        RECT 8.320 27.620 8.600 28.450 ;
        RECT 19.235 28.345 19.630 28.450 ;
        RECT 21.660 28.345 21.980 28.370 ;
        RECT 19.235 28.135 21.980 28.345 ;
        RECT 20.195 27.880 20.405 28.135 ;
        RECT 21.660 28.110 21.980 28.135 ;
        RECT 20.010 27.650 21.570 27.880 ;
        RECT 8.300 27.360 10.640 27.620 ;
        RECT 8.300 27.260 8.600 27.360 ;
        RECT 0.640 26.990 0.960 27.020 ;
        RECT 2.000 26.990 2.230 27.135 ;
        RECT 0.640 26.790 2.230 26.990 ;
        RECT 0.640 26.760 0.960 26.790 ;
        RECT 2.000 26.595 2.230 26.790 ;
        RECT 8.300 26.160 8.560 27.260 ;
        RECT 20.910 26.770 21.140 26.935 ;
        RECT 21.660 26.770 21.980 26.795 ;
        RECT 20.910 26.560 21.980 26.770 ;
        RECT 9.490 26.450 9.750 26.480 ;
        RECT 9.490 26.190 10.650 26.450 ;
        RECT 20.910 26.395 21.140 26.560 ;
        RECT 21.660 26.535 21.980 26.560 ;
        RECT 9.490 26.160 9.750 26.190 ;
        RECT -0.725 15.885 -0.375 15.915 ;
        RECT 7.020 15.885 8.020 16.020 ;
        RECT -0.725 15.535 8.020 15.885 ;
        RECT -0.725 15.505 -0.375 15.535 ;
        RECT -3.780 15.015 -3.370 15.365 ;
        RECT 7.020 15.010 8.020 15.535 ;
        RECT 16.095 15.105 26.535 15.335 ;
        RECT 2.360 14.860 15.220 15.010 ;
        RECT 2.240 14.855 15.220 14.860 ;
        RECT 16.095 14.855 16.325 15.105 ;
        RECT 2.240 14.840 16.325 14.855 ;
        RECT 1.740 14.640 16.325 14.840 ;
        RECT 1.740 14.270 1.940 14.640 ;
        RECT 2.240 14.625 16.325 14.640 ;
        RECT 2.240 14.580 15.220 14.625 ;
        RECT 2.240 14.280 4.120 14.580 ;
        RECT 1.680 14.010 2.000 14.270 ;
        RECT 2.230 14.110 4.120 14.280 ;
        RECT 2.230 14.050 3.790 14.110 ;
        RECT 8.390 13.680 8.670 14.580 ;
        RECT 26.305 14.395 26.535 15.105 ;
        RECT 23.735 14.290 26.945 14.395 ;
        RECT 23.695 14.165 26.945 14.290 ;
        RECT 23.695 14.060 23.985 14.165 ;
        RECT 23.960 13.840 24.190 13.900 ;
        RECT 25.240 13.840 25.450 14.165 ;
        RECT 8.990 13.680 11.530 13.840 ;
        RECT 8.390 13.560 11.530 13.680 ;
        RECT 23.960 13.630 25.450 13.840 ;
        RECT 8.390 13.400 9.270 13.560 ;
        RECT 23.960 13.480 24.190 13.630 ;
        RECT 1.680 13.140 2.000 13.170 ;
        RECT 2.660 13.140 2.890 13.335 ;
        RECT 1.680 12.940 2.890 13.140 ;
        RECT 1.680 12.910 2.000 12.940 ;
        RECT 2.660 12.795 2.890 12.940 ;
        RECT 8.990 12.360 9.270 13.400 ;
        RECT 23.695 13.290 23.985 13.320 ;
        RECT 24.380 13.290 25.345 13.345 ;
        RECT 23.695 13.115 25.345 13.290 ;
        RECT 23.695 13.090 23.985 13.115 ;
        RECT 25.115 13.005 25.345 13.115 ;
        RECT 26.715 13.005 26.945 14.165 ;
        RECT 29.690 13.290 34.460 13.520 ;
        RECT 29.690 13.005 29.920 13.290 ;
        RECT 34.095 13.280 34.385 13.290 ;
        RECT 25.115 12.775 29.920 13.005 ;
        RECT 10.180 12.670 10.460 12.700 ;
        RECT 10.180 12.390 11.600 12.670 ;
        RECT 29.690 12.495 29.920 12.775 ;
        RECT 34.095 12.495 34.385 12.540 ;
        RECT 10.180 12.360 10.460 12.390 ;
        RECT 29.690 12.265 34.455 12.495 ;
      LAYER met2 ;
        RECT 22.455 30.195 22.785 30.225 ;
        RECT 22.455 29.865 26.895 30.195 ;
        RECT 22.455 29.835 22.785 29.865 ;
        RECT 0.670 27.810 0.930 28.130 ;
        RECT 21.690 28.080 21.950 28.400 ;
        RECT 0.700 27.050 0.900 27.810 ;
        RECT 0.670 26.730 0.930 27.050 ;
        RECT 21.715 26.825 21.925 28.080 ;
        RECT 21.690 26.505 21.950 26.825 ;
        RECT 8.270 26.190 9.780 26.450 ;
        RECT -0.755 15.535 -0.345 15.885 ;
        RECT -3.750 15.365 -3.400 15.395 ;
        RECT -0.725 15.365 -0.375 15.535 ;
        RECT -3.750 15.015 -0.375 15.365 ;
        RECT -3.750 14.985 -3.400 15.015 ;
        RECT 1.710 13.980 1.970 14.300 ;
        RECT 1.740 13.200 1.940 13.980 ;
        RECT 1.710 12.880 1.970 13.200 ;
        RECT 8.960 12.390 10.490 12.670 ;
    END
  END VDD
  PIN down
    ANTENNAGATEAREA 2.872800 ;
    PORT
      LAYER li1 ;
        RECT 2.845 13.570 3.175 13.740 ;
        RECT 2.845 12.390 3.175 12.560 ;
        RECT 2.735 10.090 3.065 10.260 ;
        RECT 2.735 9.120 3.065 9.290 ;
        RECT 14.590 -0.105 14.760 0.225 ;
        RECT 30.140 -0.105 30.310 0.225 ;
      LAYER met1 ;
        RECT 2.865 13.760 3.155 13.770 ;
        RECT 0.640 13.550 3.170 13.760 ;
        RECT 0.640 12.515 0.850 13.550 ;
        RECT 2.865 13.540 3.155 13.550 ;
        RECT 2.865 12.515 3.155 12.590 ;
        RECT 0.640 12.305 3.195 12.515 ;
        RECT -1.240 11.600 -0.240 11.800 ;
        RECT 0.640 11.600 0.850 12.305 ;
        RECT -1.240 11.320 0.850 11.600 ;
        RECT -1.240 10.800 -0.240 11.320 ;
        RECT 0.030 4.740 0.310 11.320 ;
        RECT 0.640 10.255 0.850 11.320 ;
        RECT 2.755 10.255 3.045 10.290 ;
        RECT 0.640 10.045 3.095 10.255 ;
        RECT 0.640 9.265 0.850 10.045 ;
        RECT 2.755 9.265 3.045 9.320 ;
        RECT 0.640 9.090 3.045 9.265 ;
        RECT 0.640 9.055 3.025 9.090 ;
        RECT 3.700 4.740 3.975 4.770 ;
        RECT 7.980 4.740 8.255 4.770 ;
        RECT 0.030 4.460 2.630 4.740 ;
        RECT 3.700 4.465 7.195 4.740 ;
        RECT 7.980 4.465 18.835 4.740 ;
        RECT 3.700 4.435 3.975 4.465 ;
        RECT 7.980 4.435 8.255 4.465 ;
        RECT 14.580 1.665 14.770 1.700 ;
        RECT 18.560 1.665 18.835 4.465 ;
        RECT 14.580 1.475 30.265 1.665 ;
        RECT 14.580 0.205 14.770 1.475 ;
        RECT 18.560 1.415 18.835 1.475 ;
        RECT 30.075 0.205 30.265 1.475 ;
        RECT 14.560 -0.085 14.790 0.205 ;
        RECT 30.075 -0.035 30.340 0.205 ;
        RECT 30.110 -0.085 30.340 -0.035 ;
        RECT 14.580 -0.130 14.770 -0.085 ;
      LAYER met2 ;
        RECT 2.320 4.740 2.600 4.770 ;
        RECT 6.890 4.740 7.165 4.770 ;
        RECT 2.320 4.465 4.005 4.740 ;
        RECT 6.890 4.465 8.285 4.740 ;
        RECT 2.320 4.430 2.600 4.465 ;
        RECT 6.890 4.435 7.165 4.465 ;
    END
  END down
  OBS
      LAYER pwell ;
        RECT 56.740 43.200 58.780 43.630 ;
        RECT 56.740 36.550 57.170 43.200 ;
        RECT 58.350 36.550 58.780 43.200 ;
      LAYER nwell ;
        RECT 100.865 40.810 105.555 42.920 ;
        RECT 121.215 40.090 125.905 42.200 ;
        RECT 149.800 40.440 154.490 42.550 ;
      LAYER pwell ;
        RECT 101.745 38.020 104.745 40.030 ;
      LAYER nwell ;
        RECT 170.150 39.720 174.840 41.830 ;
      LAYER pwell ;
        RECT 121.935 37.270 124.935 39.280 ;
        RECT 150.680 37.650 153.680 39.660 ;
        RECT 170.870 36.900 173.870 38.910 ;
        RECT 56.740 36.120 58.780 36.550 ;
      LAYER nwell ;
        RECT 87.530 29.470 89.640 34.160 ;
        RECT 91.555 29.900 96.245 32.010 ;
        RECT 101.035 29.270 103.145 33.960 ;
        RECT 106.485 29.260 108.595 33.950 ;
        RECT 111.255 30.380 115.945 32.490 ;
      LAYER pwell ;
        RECT 1.350 22.820 3.390 25.240 ;
      LAYER nwell ;
        RECT 9.410 24.090 11.550 28.280 ;
        RECT 25.430 25.420 27.570 28.150 ;
      LAYER pwell ;
        RECT 87.560 25.890 89.570 28.890 ;
        RECT 92.345 27.090 95.345 29.100 ;
        RECT 101.115 26.100 103.125 29.100 ;
        RECT 106.595 25.720 108.605 28.720 ;
        RECT 112.145 27.670 115.145 29.680 ;
      LAYER nwell ;
        RECT 119.845 29.630 121.955 34.320 ;
        RECT 124.865 29.400 126.975 34.090 ;
      LAYER pwell ;
        RECT 119.925 26.360 121.935 29.360 ;
      LAYER nwell ;
        RECT 136.465 29.100 138.575 33.790 ;
        RECT 140.490 29.530 145.180 31.640 ;
      LAYER pwell ;
        RECT 124.945 26.060 126.955 29.060 ;
      LAYER nwell ;
        RECT 149.970 28.900 152.080 33.590 ;
        RECT 155.420 28.890 157.530 33.580 ;
        RECT 160.190 30.010 164.880 32.120 ;
      LAYER pwell ;
        RECT 136.495 25.520 138.505 28.520 ;
        RECT 141.280 26.720 144.280 28.730 ;
        RECT 150.050 25.730 152.060 28.730 ;
        RECT 155.530 25.350 157.540 28.350 ;
        RECT 161.080 27.300 164.080 29.310 ;
      LAYER nwell ;
        RECT 168.780 29.260 170.890 33.950 ;
        RECT 173.800 29.030 175.910 33.720 ;
      LAYER pwell ;
        RECT 168.860 25.990 170.870 28.990 ;
        RECT 173.880 25.690 175.890 28.690 ;
      LAYER nwell ;
        RECT 9.350 24.080 11.550 24.090 ;
        RECT 7.600 22.650 13.410 24.080 ;
        RECT 7.600 20.080 9.030 22.650 ;
      LAYER pwell ;
        RECT 9.480 20.160 11.520 22.580 ;
      LAYER nwell ;
        RECT 11.980 20.080 13.410 22.650 ;
        RECT 7.600 18.650 13.410 20.080 ;
        RECT 17.540 17.930 19.680 20.660 ;
      LAYER pwell ;
        RECT 1.880 8.480 3.920 10.900 ;
      LAYER nwell ;
        RECT 10.300 9.500 12.440 14.500 ;
      LAYER pwell ;
        RECT 22.820 12.480 24.860 14.900 ;
      LAYER nwell ;
        RECT 31.310 14.180 37.120 15.610 ;
      LAYER pwell ;
        RECT 116.705 15.405 118.715 18.405 ;
        RECT 121.725 15.105 123.735 18.105 ;
      LAYER nwell ;
        RECT 31.310 11.610 32.740 14.180 ;
      LAYER pwell ;
        RECT 33.220 11.700 35.260 14.120 ;
      LAYER nwell ;
        RECT 35.690 11.610 37.120 14.180 ;
        RECT 8.660 8.070 14.470 9.500 ;
        RECT 8.660 5.500 10.090 8.070 ;
      LAYER pwell ;
        RECT 10.460 5.560 12.500 7.980 ;
      LAYER nwell ;
        RECT 13.040 5.500 14.470 8.070 ;
        RECT 8.660 4.070 14.470 5.500 ;
        RECT 19.980 9.380 25.790 10.810 ;
        RECT 31.310 10.180 37.120 11.610 ;
        RECT 19.980 6.810 21.410 9.380 ;
      LAYER pwell ;
        RECT 21.920 6.870 23.960 9.290 ;
      LAYER nwell ;
        RECT 24.360 6.810 25.790 9.380 ;
        RECT 19.980 5.380 25.790 6.810 ;
        RECT 45.240 5.185 47.380 9.175 ;
        RECT 54.000 5.195 56.140 10.925 ;
        RECT 61.590 5.245 63.730 10.975 ;
        RECT 69.200 5.265 71.340 10.995 ;
        RECT 77.200 5.225 79.340 10.955 ;
        RECT 85.010 5.245 87.150 10.975 ;
        RECT 92.600 5.225 94.740 10.955 ;
        RECT 99.990 5.195 102.130 10.925 ;
        RECT 116.685 10.375 118.795 15.065 ;
        RECT 121.705 10.145 123.815 14.835 ;
      LAYER pwell ;
        RECT 128.515 14.785 131.515 16.795 ;
        RECT 135.055 15.745 137.065 18.745 ;
        RECT 140.535 15.365 142.545 18.365 ;
        RECT 148.315 15.365 151.315 17.375 ;
        RECT 154.090 15.575 156.100 18.575 ;
      LAYER nwell ;
        RECT 127.715 11.975 132.405 14.085 ;
        RECT 135.065 10.515 137.175 15.205 ;
        RECT 140.515 10.505 142.625 15.195 ;
        RECT 147.415 12.455 152.105 14.565 ;
        RECT 154.020 10.305 156.130 14.995 ;
        RECT 106.510 5.885 108.650 8.795 ;
      LAYER pwell ;
        RECT 45.280 1.845 47.320 4.265 ;
        RECT 54.060 2.485 56.100 4.905 ;
        RECT 61.650 2.535 63.690 4.955 ;
        RECT 69.260 2.555 71.300 4.975 ;
        RECT 13.950 -0.960 30.950 1.080 ;
        RECT 54.070 0.055 56.110 2.475 ;
        RECT 61.660 0.105 63.700 2.525 ;
        RECT 69.270 0.125 71.310 2.545 ;
        RECT 77.260 2.515 79.300 4.935 ;
        RECT 85.070 2.535 87.110 4.955 ;
        RECT 77.270 0.085 79.310 2.505 ;
        RECT 85.080 0.105 87.120 2.525 ;
        RECT 92.660 2.515 94.700 4.935 ;
        RECT 92.670 0.085 94.710 2.505 ;
        RECT 100.050 2.485 102.090 4.905 ;
        RECT 106.510 2.935 108.550 5.355 ;
        RECT 118.725 5.185 121.725 7.195 ;
        RECT 138.915 4.435 141.915 6.445 ;
        RECT 100.060 0.055 102.100 2.475 ;
      LAYER nwell ;
        RECT 117.755 2.265 122.445 4.375 ;
        RECT 138.105 1.545 142.795 3.655 ;
      LAYER li1 ;
        RECT 56.870 43.330 58.650 43.500 ;
        RECT 56.870 36.420 57.040 43.330 ;
        RECT 57.520 42.600 58.000 42.770 ;
        RECT 57.600 40.785 57.920 42.600 ;
        RECT 58.480 36.420 58.650 43.330 ;
        RECT 101.045 42.570 105.375 42.740 ;
        RECT 101.045 41.160 101.215 42.570 ;
        RECT 105.205 42.250 105.375 42.570 ;
        RECT 101.555 41.700 101.725 42.030 ;
        RECT 101.940 42.000 104.480 42.170 ;
        RECT 101.940 41.560 104.480 41.730 ;
        RECT 104.695 41.700 104.865 42.030 ;
        RECT 105.205 41.500 105.515 42.250 ;
        RECT 149.980 42.200 154.310 42.370 ;
        RECT 121.395 41.850 125.725 42.020 ;
        RECT 105.205 41.160 105.375 41.500 ;
        RECT 101.045 40.990 105.375 41.160 ;
        RECT 121.395 40.440 121.565 41.850 ;
        RECT 121.905 40.980 122.075 41.310 ;
        RECT 122.290 41.280 124.830 41.450 ;
        RECT 122.290 40.840 124.830 41.010 ;
        RECT 125.045 40.980 125.215 41.310 ;
        RECT 125.555 40.440 125.725 41.850 ;
        RECT 149.980 40.790 150.150 42.200 ;
        RECT 154.140 41.880 154.310 42.200 ;
        RECT 150.490 41.330 150.660 41.660 ;
        RECT 150.875 41.630 153.415 41.800 ;
        RECT 150.875 41.190 153.415 41.360 ;
        RECT 153.630 41.330 153.800 41.660 ;
        RECT 154.140 41.130 154.450 41.880 ;
        RECT 170.330 41.480 174.660 41.650 ;
        RECT 154.140 40.790 154.310 41.130 ;
        RECT 149.980 40.620 154.310 40.790 ;
        RECT 121.395 40.270 125.725 40.440 ;
        RECT 170.330 40.070 170.500 41.480 ;
        RECT 170.840 40.610 171.010 40.940 ;
        RECT 171.225 40.910 173.765 41.080 ;
        RECT 171.225 40.470 173.765 40.640 ;
        RECT 173.980 40.610 174.150 40.940 ;
        RECT 174.490 40.070 174.660 41.480 ;
        RECT 170.330 39.900 174.660 40.070 ;
        RECT 101.875 39.730 104.615 39.900 ;
        RECT 101.875 39.490 102.045 39.730 ;
        RECT 101.675 38.590 102.045 39.490 ;
        RECT 102.385 38.860 102.555 39.190 ;
        RECT 102.725 39.160 103.765 39.330 ;
        RECT 102.725 38.720 103.765 38.890 ;
        RECT 103.935 38.860 104.105 39.190 ;
        RECT 101.875 38.320 102.045 38.590 ;
        RECT 104.445 38.320 104.615 39.730 ;
        RECT 150.810 39.360 153.550 39.530 ;
        RECT 122.065 38.980 124.805 39.150 ;
        RECT 150.810 39.120 150.980 39.360 ;
        RECT 122.065 38.760 122.235 38.980 ;
        RECT 101.875 38.150 104.615 38.320 ;
        RECT 122.055 37.880 122.255 38.760 ;
        RECT 122.575 38.110 122.745 38.440 ;
        RECT 122.915 38.410 123.955 38.580 ;
        RECT 122.915 37.970 123.955 38.140 ;
        RECT 124.125 38.110 124.295 38.440 ;
        RECT 122.065 37.570 122.235 37.880 ;
        RECT 124.635 37.570 124.805 38.980 ;
        RECT 150.610 38.220 150.980 39.120 ;
        RECT 151.320 38.490 151.490 38.820 ;
        RECT 151.660 38.790 152.700 38.960 ;
        RECT 151.660 38.350 152.700 38.520 ;
        RECT 152.870 38.490 153.040 38.820 ;
        RECT 150.810 37.950 150.980 38.220 ;
        RECT 153.380 37.950 153.550 39.360 ;
        RECT 171.000 38.610 173.740 38.780 ;
        RECT 171.000 38.390 171.170 38.610 ;
        RECT 150.810 37.780 153.550 37.950 ;
        RECT 122.065 37.400 124.805 37.570 ;
        RECT 170.990 37.510 171.190 38.390 ;
        RECT 171.510 37.740 171.680 38.070 ;
        RECT 171.850 38.040 172.890 38.210 ;
        RECT 171.850 37.600 172.890 37.770 ;
        RECT 173.060 37.740 173.230 38.070 ;
        RECT 171.000 37.200 171.170 37.510 ;
        RECT 173.570 37.200 173.740 38.610 ;
        RECT 171.000 37.030 173.740 37.200 ;
        RECT 56.870 36.250 58.650 36.420 ;
        RECT 120.445 34.140 121.355 34.300 ;
        RECT 88.120 33.980 89.090 34.110 ;
        RECT 87.710 33.810 89.460 33.980 ;
        RECT 120.025 33.970 121.775 34.140 ;
        RECT -5.100 32.935 -4.930 33.265 ;
        RECT -4.715 32.780 40.325 32.950 ;
        RECT 40.540 32.935 40.710 33.265 ;
        RECT 87.710 29.820 87.880 33.810 ;
        RECT 88.420 33.300 88.750 33.470 ;
        RECT 88.280 30.545 88.450 33.085 ;
        RECT 88.720 30.545 88.890 33.085 ;
        RECT 88.420 30.160 88.750 30.330 ;
        RECT 89.290 29.820 89.460 33.810 ;
        RECT 101.635 33.780 102.575 33.820 ;
        RECT 101.215 33.610 102.965 33.780 ;
        RECT 106.995 33.770 107.965 33.910 ;
        RECT 91.735 31.660 96.065 31.830 ;
        RECT 91.735 30.250 91.905 31.660 ;
        RECT 95.895 31.400 96.065 31.660 ;
        RECT 92.245 30.790 92.415 31.120 ;
        RECT 92.630 31.090 95.170 31.260 ;
        RECT 92.630 30.650 95.170 30.820 ;
        RECT 95.385 30.790 95.555 31.120 ;
        RECT 95.895 30.550 96.130 31.400 ;
        RECT 95.895 30.250 96.065 30.550 ;
        RECT 91.735 30.080 96.065 30.250 ;
        RECT 87.710 29.650 89.460 29.820 ;
        RECT 101.215 29.620 101.385 33.610 ;
        RECT 101.925 33.100 102.255 33.270 ;
        RECT 101.785 30.345 101.955 32.885 ;
        RECT 102.225 30.345 102.395 32.885 ;
        RECT 101.925 29.960 102.255 30.130 ;
        RECT 102.795 29.620 102.965 33.610 ;
        RECT 101.215 29.450 102.965 29.620 ;
        RECT 106.665 33.600 108.415 33.770 ;
        RECT 106.665 29.610 106.835 33.600 ;
        RECT 107.375 33.090 107.705 33.260 ;
        RECT 107.235 30.335 107.405 32.875 ;
        RECT 107.675 30.335 107.845 32.875 ;
        RECT 107.375 29.950 107.705 30.120 ;
        RECT 108.245 29.610 108.415 33.600 ;
        RECT 111.435 32.140 115.765 32.310 ;
        RECT 111.435 30.730 111.605 32.140 ;
        RECT 115.595 32.000 115.765 32.140 ;
        RECT 111.945 31.270 112.115 31.600 ;
        RECT 112.330 31.570 114.870 31.740 ;
        RECT 112.330 31.130 114.870 31.300 ;
        RECT 115.085 31.270 115.255 31.600 ;
        RECT 115.595 30.890 115.875 32.000 ;
        RECT 115.595 30.730 115.765 30.890 ;
        RECT 111.435 30.560 115.765 30.730 ;
        RECT 120.025 29.980 120.195 33.970 ;
        RECT 120.445 33.960 121.355 33.970 ;
        RECT 120.735 33.460 121.065 33.630 ;
        RECT 120.595 30.705 120.765 33.245 ;
        RECT 121.035 30.705 121.205 33.245 ;
        RECT 120.735 30.320 121.065 30.490 ;
        RECT 121.605 29.980 121.775 33.970 ;
        RECT 125.450 33.910 126.420 34.060 ;
        RECT 120.025 29.810 121.775 29.980 ;
        RECT 125.045 33.740 126.795 33.910 ;
        RECT 169.380 33.770 170.290 33.930 ;
        RECT 106.665 29.440 108.415 29.610 ;
        RECT 125.045 29.750 125.215 33.740 ;
        RECT 125.755 33.230 126.085 33.400 ;
        RECT 125.615 30.475 125.785 33.015 ;
        RECT 126.055 30.475 126.225 33.015 ;
        RECT 125.755 30.090 126.085 30.260 ;
        RECT 126.625 29.750 126.795 33.740 ;
        RECT 137.055 33.610 138.025 33.740 ;
        RECT 125.045 29.580 126.795 29.750 ;
        RECT 136.645 33.440 138.395 33.610 ;
        RECT 168.960 33.600 170.710 33.770 ;
        RECT 112.275 29.380 115.015 29.550 ;
        RECT 112.275 29.220 112.445 29.380 ;
        RECT 92.475 28.800 95.215 28.970 ;
        RECT 87.690 28.590 89.440 28.760 ;
        RECT 9.590 27.930 11.370 28.100 ;
        RECT 2.500 26.575 2.670 27.155 ;
        RECT 9.590 25.900 9.760 27.930 ;
        RECT 10.160 26.625 10.330 27.205 ;
        RECT 10.630 26.625 10.800 27.205 ;
        RECT 11.200 25.900 11.370 27.930 ;
        RECT 25.610 27.800 27.390 27.970 ;
        RECT 20.625 27.170 20.955 27.340 ;
        RECT 20.470 26.375 20.640 26.955 ;
        RECT 20.625 25.990 20.955 26.160 ;
        RECT 9.590 25.730 11.370 25.900 ;
        RECT 25.610 25.770 25.780 27.800 ;
        RECT 26.335 27.290 26.665 27.460 ;
        RECT 26.180 26.495 26.350 27.075 ;
        RECT 26.335 26.110 26.665 26.280 ;
        RECT 27.220 25.770 27.390 27.800 ;
        RECT 87.690 26.190 87.860 28.590 ;
        RECT 88.400 28.080 88.730 28.250 ;
        RECT 88.260 26.870 88.430 27.910 ;
        RECT 88.700 26.870 88.870 27.910 ;
        RECT 88.400 26.530 88.730 26.700 ;
        RECT 89.270 26.190 89.440 28.590 ;
        RECT 92.475 28.560 92.645 28.800 ;
        RECT 92.390 27.700 92.645 28.560 ;
        RECT 92.985 27.930 93.155 28.260 ;
        RECT 93.325 28.230 94.365 28.400 ;
        RECT 93.325 27.790 94.365 27.960 ;
        RECT 94.535 27.930 94.705 28.260 ;
        RECT 92.475 27.390 92.645 27.700 ;
        RECT 95.045 27.390 95.215 28.800 ;
        RECT 92.475 27.220 95.215 27.390 ;
        RECT 101.245 28.800 102.995 28.970 ;
        RECT 101.245 26.400 101.415 28.800 ;
        RECT 101.955 28.290 102.285 28.460 ;
        RECT 101.815 27.080 101.985 28.120 ;
        RECT 102.255 27.080 102.425 28.120 ;
        RECT 101.955 26.740 102.285 26.910 ;
        RECT 102.825 26.400 102.995 28.800 ;
        RECT 101.245 26.230 102.995 26.400 ;
        RECT 106.725 28.420 108.475 28.590 ;
        RECT 87.690 26.020 89.440 26.190 ;
        RECT 101.685 26.160 102.555 26.230 ;
        RECT 106.725 26.020 106.895 28.420 ;
        RECT 107.435 27.910 107.765 28.080 ;
        RECT 107.295 26.700 107.465 27.740 ;
        RECT 107.735 26.700 107.905 27.740 ;
        RECT 107.435 26.360 107.765 26.530 ;
        RECT 108.305 26.020 108.475 28.420 ;
        RECT 112.215 28.250 112.445 29.220 ;
        RECT 112.785 28.510 112.955 28.840 ;
        RECT 113.125 28.810 114.165 28.980 ;
        RECT 113.125 28.370 114.165 28.540 ;
        RECT 114.335 28.510 114.505 28.840 ;
        RECT 112.275 27.970 112.445 28.250 ;
        RECT 114.845 27.970 115.015 29.380 ;
        RECT 136.645 29.450 136.815 33.440 ;
        RECT 137.355 32.930 137.685 33.100 ;
        RECT 137.215 30.175 137.385 32.715 ;
        RECT 137.655 30.175 137.825 32.715 ;
        RECT 137.355 29.790 137.685 29.960 ;
        RECT 138.225 29.450 138.395 33.440 ;
        RECT 150.570 33.410 151.510 33.450 ;
        RECT 150.150 33.240 151.900 33.410 ;
        RECT 155.930 33.400 156.900 33.540 ;
        RECT 140.670 31.290 145.000 31.460 ;
        RECT 140.670 29.880 140.840 31.290 ;
        RECT 144.830 31.030 145.000 31.290 ;
        RECT 141.180 30.420 141.350 30.750 ;
        RECT 141.565 30.720 144.105 30.890 ;
        RECT 141.565 30.280 144.105 30.450 ;
        RECT 144.320 30.420 144.490 30.750 ;
        RECT 144.830 30.180 145.065 31.030 ;
        RECT 144.830 29.880 145.000 30.180 ;
        RECT 140.670 29.710 145.000 29.880 ;
        RECT 136.645 29.280 138.395 29.450 ;
        RECT 150.150 29.250 150.320 33.240 ;
        RECT 150.860 32.730 151.190 32.900 ;
        RECT 150.720 29.975 150.890 32.515 ;
        RECT 151.160 29.975 151.330 32.515 ;
        RECT 150.860 29.590 151.190 29.760 ;
        RECT 151.730 29.250 151.900 33.240 ;
        RECT 112.275 27.800 115.015 27.970 ;
        RECT 120.055 29.060 121.805 29.230 ;
        RECT 150.150 29.080 151.900 29.250 ;
        RECT 155.600 33.230 157.350 33.400 ;
        RECT 155.600 29.240 155.770 33.230 ;
        RECT 156.310 32.720 156.640 32.890 ;
        RECT 156.170 29.965 156.340 32.505 ;
        RECT 156.610 29.965 156.780 32.505 ;
        RECT 156.310 29.580 156.640 29.750 ;
        RECT 157.180 29.240 157.350 33.230 ;
        RECT 160.370 31.770 164.700 31.940 ;
        RECT 160.370 30.360 160.540 31.770 ;
        RECT 164.530 31.630 164.700 31.770 ;
        RECT 160.880 30.900 161.050 31.230 ;
        RECT 161.265 31.200 163.805 31.370 ;
        RECT 161.265 30.760 163.805 30.930 ;
        RECT 164.020 30.900 164.190 31.230 ;
        RECT 164.530 30.520 164.810 31.630 ;
        RECT 164.530 30.360 164.700 30.520 ;
        RECT 160.370 30.190 164.700 30.360 ;
        RECT 168.960 29.610 169.130 33.600 ;
        RECT 169.380 33.590 170.290 33.600 ;
        RECT 169.670 33.090 170.000 33.260 ;
        RECT 169.530 30.335 169.700 32.875 ;
        RECT 169.970 30.335 170.140 32.875 ;
        RECT 169.670 29.950 170.000 30.120 ;
        RECT 170.540 29.610 170.710 33.600 ;
        RECT 174.385 33.540 175.355 33.690 ;
        RECT 168.960 29.440 170.710 29.610 ;
        RECT 173.980 33.370 175.730 33.540 ;
        RECT 155.600 29.070 157.350 29.240 ;
        RECT 173.980 29.380 174.150 33.370 ;
        RECT 174.690 32.860 175.020 33.030 ;
        RECT 174.550 30.105 174.720 32.645 ;
        RECT 174.990 30.105 175.160 32.645 ;
        RECT 174.690 29.720 175.020 29.890 ;
        RECT 175.560 29.380 175.730 33.370 ;
        RECT 173.980 29.210 175.730 29.380 ;
        RECT 120.055 26.660 120.225 29.060 ;
        RECT 120.765 28.550 121.095 28.720 ;
        RECT 120.625 27.340 120.795 28.380 ;
        RECT 121.065 27.340 121.235 28.380 ;
        RECT 120.765 27.000 121.095 27.170 ;
        RECT 121.635 26.660 121.805 29.060 ;
        RECT 161.210 29.010 163.950 29.180 ;
        RECT 120.055 26.490 121.805 26.660 ;
        RECT 125.075 28.760 126.825 28.930 ;
        RECT 161.210 28.850 161.380 29.010 ;
        RECT 120.510 26.410 121.340 26.490 ;
        RECT 125.075 26.360 125.245 28.760 ;
        RECT 125.785 28.250 126.115 28.420 ;
        RECT 125.645 27.040 125.815 28.080 ;
        RECT 126.085 27.040 126.255 28.080 ;
        RECT 125.785 26.700 126.115 26.870 ;
        RECT 126.655 26.360 126.825 28.760 ;
        RECT 141.410 28.430 144.150 28.600 ;
        RECT 125.075 26.190 126.825 26.360 ;
        RECT 136.625 28.220 138.375 28.390 ;
        RECT 125.510 26.070 126.370 26.190 ;
        RECT 88.140 25.960 88.990 26.020 ;
        RECT 106.725 25.850 108.475 26.020 ;
        RECT 25.610 25.600 27.390 25.770 ;
        RECT 107.050 25.740 108.140 25.850 ;
        RECT 136.625 25.820 136.795 28.220 ;
        RECT 137.335 27.710 137.665 27.880 ;
        RECT 137.195 26.500 137.365 27.540 ;
        RECT 137.635 26.500 137.805 27.540 ;
        RECT 137.335 26.160 137.665 26.330 ;
        RECT 138.205 25.820 138.375 28.220 ;
        RECT 141.410 28.190 141.580 28.430 ;
        RECT 141.325 27.330 141.580 28.190 ;
        RECT 141.920 27.560 142.090 27.890 ;
        RECT 142.260 27.860 143.300 28.030 ;
        RECT 142.260 27.420 143.300 27.590 ;
        RECT 143.470 27.560 143.640 27.890 ;
        RECT 141.410 27.020 141.580 27.330 ;
        RECT 143.980 27.020 144.150 28.430 ;
        RECT 141.410 26.850 144.150 27.020 ;
        RECT 150.180 28.430 151.930 28.600 ;
        RECT 150.180 26.030 150.350 28.430 ;
        RECT 150.890 27.920 151.220 28.090 ;
        RECT 150.750 26.710 150.920 27.750 ;
        RECT 151.190 26.710 151.360 27.750 ;
        RECT 150.890 26.370 151.220 26.540 ;
        RECT 151.760 26.030 151.930 28.430 ;
        RECT 150.180 25.860 151.930 26.030 ;
        RECT 155.660 28.050 157.410 28.220 ;
        RECT 136.625 25.650 138.375 25.820 ;
        RECT 150.620 25.790 151.490 25.860 ;
        RECT 155.660 25.650 155.830 28.050 ;
        RECT 156.370 27.540 156.700 27.710 ;
        RECT 156.230 26.330 156.400 27.370 ;
        RECT 156.670 26.330 156.840 27.370 ;
        RECT 156.370 25.990 156.700 26.160 ;
        RECT 157.240 25.650 157.410 28.050 ;
        RECT 161.150 27.880 161.380 28.850 ;
        RECT 161.720 28.140 161.890 28.470 ;
        RECT 162.060 28.440 163.100 28.610 ;
        RECT 162.060 28.000 163.100 28.170 ;
        RECT 163.270 28.140 163.440 28.470 ;
        RECT 161.210 27.600 161.380 27.880 ;
        RECT 163.780 27.600 163.950 29.010 ;
        RECT 161.210 27.430 163.950 27.600 ;
        RECT 168.990 28.690 170.740 28.860 ;
        RECT 168.990 26.290 169.160 28.690 ;
        RECT 169.700 28.180 170.030 28.350 ;
        RECT 169.560 26.970 169.730 28.010 ;
        RECT 170.000 26.970 170.170 28.010 ;
        RECT 169.700 26.630 170.030 26.800 ;
        RECT 170.570 26.290 170.740 28.690 ;
        RECT 168.990 26.120 170.740 26.290 ;
        RECT 174.010 28.390 175.760 28.560 ;
        RECT 169.445 26.040 170.275 26.120 ;
        RECT 174.010 25.990 174.180 28.390 ;
        RECT 174.720 27.880 175.050 28.050 ;
        RECT 174.580 26.670 174.750 27.710 ;
        RECT 175.020 26.670 175.190 27.710 ;
        RECT 174.720 26.330 175.050 26.500 ;
        RECT 175.590 25.990 175.760 28.390 ;
        RECT 174.010 25.820 175.760 25.990 ;
        RECT 174.445 25.700 175.305 25.820 ;
        RECT 137.075 25.590 137.925 25.650 ;
        RECT 155.660 25.480 157.410 25.650 ;
        RECT 155.985 25.370 157.075 25.480 ;
        RECT 1.480 24.940 3.260 25.110 ;
        RECT 1.480 23.120 1.650 24.940 ;
        RECT 2.050 23.800 2.220 24.260 ;
        RECT 2.520 23.800 2.690 24.260 ;
        RECT 3.090 23.120 3.260 24.940 ;
        RECT 1.480 22.950 3.260 23.120 ;
        RECT 7.885 23.625 13.125 23.795 ;
        RECT 7.885 19.105 8.055 23.625 ;
        RECT 9.610 22.280 11.390 22.450 ;
        RECT 9.610 20.460 9.780 22.280 ;
        RECT 10.335 21.770 10.665 21.940 ;
        RECT 10.180 21.140 10.350 21.600 ;
        RECT 10.650 21.140 10.820 21.600 ;
        RECT 10.335 20.800 10.665 20.970 ;
        RECT 11.220 20.460 11.390 22.280 ;
        RECT 9.610 20.290 11.390 20.460 ;
        RECT 12.955 19.105 13.125 23.625 ;
        RECT 7.885 18.935 13.125 19.105 ;
        RECT 17.720 20.310 19.500 20.480 ;
        RECT 17.720 18.280 17.890 20.310 ;
        RECT 18.290 19.005 18.460 19.585 ;
        RECT 18.760 19.005 18.930 19.585 ;
        RECT 19.330 18.280 19.500 20.310 ;
        RECT 135.520 18.615 136.610 18.725 ;
        RECT 135.185 18.445 136.935 18.615 ;
        RECT 154.670 18.445 155.520 18.505 ;
        RECT 17.720 18.110 19.500 18.280 ;
        RECT 117.290 18.275 118.150 18.395 ;
        RECT 116.835 18.105 118.585 18.275 ;
        RECT 116.835 15.705 117.005 18.105 ;
        RECT 117.545 17.595 117.875 17.765 ;
        RECT 117.405 16.385 117.575 17.425 ;
        RECT 117.845 16.385 118.015 17.425 ;
        RECT 117.545 16.045 117.875 16.215 ;
        RECT 118.415 15.705 118.585 18.105 ;
        RECT 122.320 17.975 123.150 18.055 ;
        RECT 116.835 15.535 118.585 15.705 ;
        RECT 121.855 17.805 123.605 17.975 ;
        RECT 121.855 15.405 122.025 17.805 ;
        RECT 122.565 17.295 122.895 17.465 ;
        RECT 122.425 16.085 122.595 17.125 ;
        RECT 122.865 16.085 123.035 17.125 ;
        RECT 122.565 15.745 122.895 15.915 ;
        RECT 123.435 15.405 123.605 17.805 ;
        RECT 31.595 15.155 36.835 15.325 ;
        RECT 121.855 15.235 123.605 15.405 ;
        RECT 128.645 16.495 131.385 16.665 ;
        RECT 22.950 14.600 24.730 14.770 ;
        RECT 10.480 14.150 12.260 14.320 ;
        RECT 3.160 12.775 3.330 13.355 ;
        RECT 10.480 12.120 10.650 14.150 ;
        RECT 11.050 12.845 11.220 13.425 ;
        RECT 11.520 12.845 11.690 13.425 ;
        RECT 12.090 12.120 12.260 14.150 ;
        RECT 22.950 12.780 23.120 14.600 ;
        RECT 23.520 13.460 23.690 13.920 ;
        RECT 24.560 12.780 24.730 14.600 ;
        RECT 22.950 12.610 24.730 12.780 ;
        RECT 10.480 11.950 12.260 12.120 ;
        RECT 2.010 10.600 3.790 10.770 ;
        RECT 2.010 8.780 2.180 10.600 ;
        RECT 2.580 9.460 2.750 9.920 ;
        RECT 3.050 9.460 3.220 9.920 ;
        RECT 3.620 8.780 3.790 10.600 ;
        RECT 31.595 10.635 31.765 15.155 ;
        RECT 33.350 13.820 35.130 13.990 ;
        RECT 33.350 12.000 33.520 13.820 ;
        RECT 34.390 12.680 34.560 13.140 ;
        RECT 34.960 12.000 35.130 13.820 ;
        RECT 33.350 11.830 35.130 12.000 ;
        RECT 36.665 10.635 36.835 15.155 ;
        RECT 128.645 15.085 128.815 16.495 ;
        RECT 131.215 16.215 131.385 16.495 ;
        RECT 129.155 15.625 129.325 15.955 ;
        RECT 129.495 15.925 130.535 16.095 ;
        RECT 129.495 15.485 130.535 15.655 ;
        RECT 130.705 15.625 130.875 15.955 ;
        RECT 131.215 15.245 131.445 16.215 ;
        RECT 135.185 16.045 135.355 18.445 ;
        RECT 135.895 17.935 136.225 18.105 ;
        RECT 135.755 16.725 135.925 17.765 ;
        RECT 136.195 16.725 136.365 17.765 ;
        RECT 135.895 16.385 136.225 16.555 ;
        RECT 136.765 16.045 136.935 18.445 ;
        RECT 141.105 18.235 141.975 18.305 ;
        RECT 154.220 18.275 155.970 18.445 ;
        RECT 135.185 15.875 136.935 16.045 ;
        RECT 140.665 18.065 142.415 18.235 ;
        RECT 140.665 15.665 140.835 18.065 ;
        RECT 141.375 17.555 141.705 17.725 ;
        RECT 141.235 16.345 141.405 17.385 ;
        RECT 141.675 16.345 141.845 17.385 ;
        RECT 141.375 16.005 141.705 16.175 ;
        RECT 142.245 15.665 142.415 18.065 ;
        RECT 140.665 15.495 142.415 15.665 ;
        RECT 148.445 17.075 151.185 17.245 ;
        RECT 148.445 15.665 148.615 17.075 ;
        RECT 151.015 16.765 151.185 17.075 ;
        RECT 148.955 16.205 149.125 16.535 ;
        RECT 149.295 16.505 150.335 16.675 ;
        RECT 149.295 16.065 150.335 16.235 ;
        RECT 150.505 16.205 150.675 16.535 ;
        RECT 151.015 15.905 151.270 16.765 ;
        RECT 151.015 15.665 151.185 15.905 ;
        RECT 154.220 15.875 154.390 18.275 ;
        RECT 154.930 17.765 155.260 17.935 ;
        RECT 154.790 16.555 154.960 17.595 ;
        RECT 155.230 16.555 155.400 17.595 ;
        RECT 154.930 16.215 155.260 16.385 ;
        RECT 155.800 15.875 155.970 18.275 ;
        RECT 154.220 15.705 155.970 15.875 ;
        RECT 148.445 15.495 151.185 15.665 ;
        RECT 131.215 15.085 131.385 15.245 ;
        RECT 128.645 14.915 131.385 15.085 ;
        RECT 116.865 14.715 118.615 14.885 ;
        RECT 54.560 10.745 55.550 10.885 ;
        RECT 62.150 10.795 63.140 10.935 ;
        RECT 69.760 10.815 70.750 10.955 ;
        RECT 20.265 10.355 25.505 10.525 ;
        RECT 31.595 10.465 36.835 10.635 ;
        RECT 54.180 10.575 55.960 10.745 ;
        RECT 2.010 8.610 3.790 8.780 ;
        RECT 8.945 9.045 14.185 9.215 ;
        RECT 8.945 4.525 9.115 9.045 ;
        RECT 10.590 7.680 12.370 7.850 ;
        RECT 10.590 5.860 10.760 7.680 ;
        RECT 11.315 7.170 11.645 7.340 ;
        RECT 11.160 6.540 11.330 7.000 ;
        RECT 11.630 6.540 11.800 7.000 ;
        RECT 11.315 6.200 11.645 6.370 ;
        RECT 12.200 5.860 12.370 7.680 ;
        RECT 10.590 5.690 12.370 5.860 ;
        RECT 14.015 4.525 14.185 9.045 ;
        RECT 20.265 5.835 20.435 10.355 ;
        RECT 22.050 8.990 23.830 9.160 ;
        RECT 22.050 7.170 22.220 8.990 ;
        RECT 22.775 8.480 23.105 8.650 ;
        RECT 22.620 7.850 22.790 8.310 ;
        RECT 23.090 7.850 23.260 8.310 ;
        RECT 22.775 7.510 23.105 7.680 ;
        RECT 23.660 7.170 23.830 8.990 ;
        RECT 22.050 7.000 23.830 7.170 ;
        RECT 25.335 5.835 25.505 10.355 ;
        RECT 20.265 5.665 25.505 5.835 ;
        RECT 45.420 8.825 47.200 8.995 ;
        RECT 45.420 5.535 45.590 8.825 ;
        RECT 46.145 8.315 46.475 8.485 ;
        RECT 45.990 6.260 46.160 8.100 ;
        RECT 46.460 6.260 46.630 8.100 ;
        RECT 46.145 5.875 46.475 6.045 ;
        RECT 47.030 5.535 47.200 8.825 ;
        RECT 54.180 8.365 54.350 10.575 ;
        RECT 54.905 10.065 55.235 10.235 ;
        RECT 54.750 9.090 54.920 9.850 ;
        RECT 55.220 9.090 55.390 9.850 ;
        RECT 54.905 8.705 55.235 8.875 ;
        RECT 55.790 8.365 55.960 10.575 ;
        RECT 54.180 8.195 55.960 8.365 ;
        RECT 61.770 10.625 63.550 10.795 ;
        RECT 61.770 8.415 61.940 10.625 ;
        RECT 62.495 10.115 62.825 10.285 ;
        RECT 62.340 9.140 62.510 9.900 ;
        RECT 62.810 9.140 62.980 9.900 ;
        RECT 62.495 8.755 62.825 8.925 ;
        RECT 63.380 8.415 63.550 10.625 ;
        RECT 61.770 8.245 63.550 8.415 ;
        RECT 69.380 10.645 71.160 10.815 ;
        RECT 77.760 10.775 78.750 10.915 ;
        RECT 85.570 10.795 86.560 10.935 ;
        RECT 69.380 8.435 69.550 10.645 ;
        RECT 70.105 10.135 70.435 10.305 ;
        RECT 69.950 9.160 70.120 9.920 ;
        RECT 70.420 9.160 70.590 9.920 ;
        RECT 70.105 8.775 70.435 8.945 ;
        RECT 70.990 8.435 71.160 10.645 ;
        RECT 69.380 8.265 71.160 8.435 ;
        RECT 77.380 10.605 79.160 10.775 ;
        RECT 77.380 8.395 77.550 10.605 ;
        RECT 78.105 10.095 78.435 10.265 ;
        RECT 77.950 9.120 78.120 9.880 ;
        RECT 78.420 9.120 78.590 9.880 ;
        RECT 78.105 8.735 78.435 8.905 ;
        RECT 78.990 8.395 79.160 10.605 ;
        RECT 77.380 8.225 79.160 8.395 ;
        RECT 85.190 10.625 86.970 10.795 ;
        RECT 93.160 10.775 94.150 10.915 ;
        RECT 85.190 8.415 85.360 10.625 ;
        RECT 85.915 10.115 86.245 10.285 ;
        RECT 85.760 9.140 85.930 9.900 ;
        RECT 86.230 9.140 86.400 9.900 ;
        RECT 85.915 8.755 86.245 8.925 ;
        RECT 86.800 8.415 86.970 10.625 ;
        RECT 85.190 8.245 86.970 8.415 ;
        RECT 92.780 10.605 94.560 10.775 ;
        RECT 100.550 10.745 101.540 10.885 ;
        RECT 92.780 8.395 92.950 10.605 ;
        RECT 93.505 10.095 93.835 10.265 ;
        RECT 93.350 9.120 93.520 9.880 ;
        RECT 93.820 9.120 93.990 9.880 ;
        RECT 93.505 8.735 93.835 8.905 ;
        RECT 94.390 8.395 94.560 10.605 ;
        RECT 92.780 8.225 94.560 8.395 ;
        RECT 100.170 10.575 101.950 10.745 ;
        RECT 100.170 8.365 100.340 10.575 ;
        RECT 100.895 10.065 101.225 10.235 ;
        RECT 100.740 9.090 100.910 9.850 ;
        RECT 101.210 9.090 101.380 9.850 ;
        RECT 100.895 8.705 101.225 8.875 ;
        RECT 101.780 8.365 101.950 10.575 ;
        RECT 116.865 10.725 117.035 14.715 ;
        RECT 117.575 14.205 117.905 14.375 ;
        RECT 117.435 11.450 117.605 13.990 ;
        RECT 117.875 11.450 118.045 13.990 ;
        RECT 117.575 11.065 117.905 11.235 ;
        RECT 118.445 10.725 118.615 14.715 ;
        RECT 135.245 14.855 136.995 15.025 ;
        RECT 116.865 10.555 118.615 10.725 ;
        RECT 121.885 14.485 123.635 14.655 ;
        RECT 117.240 10.405 118.210 10.555 ;
        RECT 121.885 10.495 122.055 14.485 ;
        RECT 122.595 13.975 122.925 14.145 ;
        RECT 122.455 11.220 122.625 13.760 ;
        RECT 122.895 11.220 123.065 13.760 ;
        RECT 122.595 10.835 122.925 11.005 ;
        RECT 122.305 10.495 123.215 10.505 ;
        RECT 123.465 10.495 123.635 14.485 ;
        RECT 127.895 13.735 132.225 13.905 ;
        RECT 127.895 13.575 128.065 13.735 ;
        RECT 127.785 12.465 128.065 13.575 ;
        RECT 128.405 12.865 128.575 13.195 ;
        RECT 128.790 13.165 131.330 13.335 ;
        RECT 128.790 12.725 131.330 12.895 ;
        RECT 131.545 12.865 131.715 13.195 ;
        RECT 127.895 12.325 128.065 12.465 ;
        RECT 132.055 12.325 132.225 13.735 ;
        RECT 127.895 12.155 132.225 12.325 ;
        RECT 135.245 10.865 135.415 14.855 ;
        RECT 135.955 14.345 136.285 14.515 ;
        RECT 135.815 11.590 135.985 14.130 ;
        RECT 136.255 11.590 136.425 14.130 ;
        RECT 135.955 11.205 136.285 11.375 ;
        RECT 136.825 10.865 136.995 14.855 ;
        RECT 135.245 10.695 136.995 10.865 ;
        RECT 140.695 14.845 142.445 15.015 ;
        RECT 140.695 10.855 140.865 14.845 ;
        RECT 141.405 14.335 141.735 14.505 ;
        RECT 141.265 11.580 141.435 14.120 ;
        RECT 141.705 11.580 141.875 14.120 ;
        RECT 141.405 11.195 141.735 11.365 ;
        RECT 142.275 10.855 142.445 14.845 ;
        RECT 154.200 14.645 155.950 14.815 ;
        RECT 147.595 14.215 151.925 14.385 ;
        RECT 147.595 13.915 147.765 14.215 ;
        RECT 147.530 13.065 147.765 13.915 ;
        RECT 148.105 13.345 148.275 13.675 ;
        RECT 148.490 13.645 151.030 13.815 ;
        RECT 148.490 13.205 151.030 13.375 ;
        RECT 151.245 13.345 151.415 13.675 ;
        RECT 147.595 12.805 147.765 13.065 ;
        RECT 151.755 12.805 151.925 14.215 ;
        RECT 147.595 12.635 151.925 12.805 ;
        RECT 135.695 10.555 136.665 10.695 ;
        RECT 140.695 10.685 142.445 10.855 ;
        RECT 141.085 10.645 142.025 10.685 ;
        RECT 154.200 10.655 154.370 14.645 ;
        RECT 154.910 14.135 155.240 14.305 ;
        RECT 154.770 11.380 154.940 13.920 ;
        RECT 155.210 11.380 155.380 13.920 ;
        RECT 154.910 10.995 155.240 11.165 ;
        RECT 155.780 10.655 155.950 14.645 ;
        RECT 121.885 10.325 123.635 10.495 ;
        RECT 154.200 10.485 155.950 10.655 ;
        RECT 154.570 10.355 155.540 10.485 ;
        RECT 122.305 10.165 123.215 10.325 ;
        RECT 107.180 8.615 108.020 8.695 ;
        RECT 100.170 8.195 101.950 8.365 ;
        RECT 106.690 8.445 108.470 8.615 ;
        RECT 45.420 5.365 47.200 5.535 ;
        RECT 54.180 7.755 55.960 7.925 ;
        RECT 54.180 5.545 54.350 7.755 ;
        RECT 54.905 7.245 55.235 7.415 ;
        RECT 54.750 6.270 54.920 7.030 ;
        RECT 55.220 6.270 55.390 7.030 ;
        RECT 54.905 5.885 55.235 6.055 ;
        RECT 55.790 5.545 55.960 7.755 ;
        RECT 54.180 5.375 55.960 5.545 ;
        RECT 61.770 7.805 63.550 7.975 ;
        RECT 61.770 5.595 61.940 7.805 ;
        RECT 62.495 7.295 62.825 7.465 ;
        RECT 62.340 6.320 62.510 7.080 ;
        RECT 62.810 6.320 62.980 7.080 ;
        RECT 62.495 5.935 62.825 6.105 ;
        RECT 63.380 5.595 63.550 7.805 ;
        RECT 61.770 5.425 63.550 5.595 ;
        RECT 69.380 7.825 71.160 7.995 ;
        RECT 69.380 5.615 69.550 7.825 ;
        RECT 70.105 7.315 70.435 7.485 ;
        RECT 69.950 6.340 70.120 7.100 ;
        RECT 70.420 6.340 70.590 7.100 ;
        RECT 70.105 5.955 70.435 6.125 ;
        RECT 70.990 5.615 71.160 7.825 ;
        RECT 69.380 5.445 71.160 5.615 ;
        RECT 77.380 7.785 79.160 7.955 ;
        RECT 77.380 5.575 77.550 7.785 ;
        RECT 78.105 7.275 78.435 7.445 ;
        RECT 77.950 6.300 78.120 7.060 ;
        RECT 78.420 6.300 78.590 7.060 ;
        RECT 78.105 5.915 78.435 6.085 ;
        RECT 78.990 5.575 79.160 7.785 ;
        RECT 77.380 5.405 79.160 5.575 ;
        RECT 85.190 7.805 86.970 7.975 ;
        RECT 85.190 5.595 85.360 7.805 ;
        RECT 85.915 7.295 86.245 7.465 ;
        RECT 85.760 6.320 85.930 7.080 ;
        RECT 86.230 6.320 86.400 7.080 ;
        RECT 85.915 5.935 86.245 6.105 ;
        RECT 86.800 5.595 86.970 7.805 ;
        RECT 85.190 5.425 86.970 5.595 ;
        RECT 92.780 7.785 94.560 7.955 ;
        RECT 92.780 5.575 92.950 7.785 ;
        RECT 93.505 7.275 93.835 7.445 ;
        RECT 93.350 6.300 93.520 7.060 ;
        RECT 93.820 6.300 93.990 7.060 ;
        RECT 93.505 5.915 93.835 6.085 ;
        RECT 94.390 5.575 94.560 7.785 ;
        RECT 92.780 5.405 94.560 5.575 ;
        RECT 100.170 7.755 101.950 7.925 ;
        RECT 100.170 5.545 100.340 7.755 ;
        RECT 100.895 7.245 101.225 7.415 ;
        RECT 100.740 6.270 100.910 7.030 ;
        RECT 101.210 6.270 101.380 7.030 ;
        RECT 100.895 5.885 101.225 6.055 ;
        RECT 101.780 5.545 101.950 7.755 ;
        RECT 106.690 6.235 106.860 8.445 ;
        RECT 107.415 7.935 107.745 8.105 ;
        RECT 107.260 6.960 107.430 7.720 ;
        RECT 107.730 6.960 107.900 7.720 ;
        RECT 107.415 6.575 107.745 6.745 ;
        RECT 108.300 6.235 108.470 8.445 ;
        RECT 106.690 6.065 108.470 6.235 ;
        RECT 118.855 6.895 121.595 7.065 ;
        RECT 100.170 5.375 101.950 5.545 ;
        RECT 118.855 5.485 119.025 6.895 ;
        RECT 121.425 6.585 121.595 6.895 ;
        RECT 119.365 6.025 119.535 6.355 ;
        RECT 119.705 6.325 120.745 6.495 ;
        RECT 119.705 5.885 120.745 6.055 ;
        RECT 120.915 6.025 121.085 6.355 ;
        RECT 121.405 5.705 121.605 6.585 ;
        RECT 139.045 6.145 141.785 6.315 ;
        RECT 121.425 5.485 121.595 5.705 ;
        RECT 118.855 5.315 121.595 5.485 ;
        RECT 106.640 5.055 108.420 5.225 ;
        RECT 8.945 4.355 14.185 4.525 ;
        RECT 54.190 4.605 55.970 4.775 ;
        RECT 45.410 3.965 47.190 4.135 ;
        RECT 45.410 2.145 45.580 3.965 ;
        RECT 46.135 3.455 46.465 3.625 ;
        RECT 45.980 2.825 46.150 3.285 ;
        RECT 46.450 2.825 46.620 3.285 ;
        RECT 46.135 2.485 46.465 2.655 ;
        RECT 47.020 2.145 47.190 3.965 ;
        RECT 54.190 2.785 54.360 4.605 ;
        RECT 54.915 4.095 55.245 4.265 ;
        RECT 54.760 3.465 54.930 3.925 ;
        RECT 55.230 3.465 55.400 3.925 ;
        RECT 54.915 3.125 55.245 3.295 ;
        RECT 55.800 2.785 55.970 4.605 ;
        RECT 54.190 2.615 55.970 2.785 ;
        RECT 61.780 4.655 63.560 4.825 ;
        RECT 61.780 2.835 61.950 4.655 ;
        RECT 62.505 4.145 62.835 4.315 ;
        RECT 62.350 3.515 62.520 3.975 ;
        RECT 62.820 3.515 62.990 3.975 ;
        RECT 62.505 3.175 62.835 3.345 ;
        RECT 63.390 2.835 63.560 4.655 ;
        RECT 61.780 2.665 63.560 2.835 ;
        RECT 69.390 4.675 71.170 4.845 ;
        RECT 69.390 2.855 69.560 4.675 ;
        RECT 70.115 4.165 70.445 4.335 ;
        RECT 69.960 3.535 70.130 3.995 ;
        RECT 70.430 3.535 70.600 3.995 ;
        RECT 70.115 3.195 70.445 3.365 ;
        RECT 71.000 2.855 71.170 4.675 ;
        RECT 69.390 2.685 71.170 2.855 ;
        RECT 77.390 4.635 79.170 4.805 ;
        RECT 77.390 2.815 77.560 4.635 ;
        RECT 78.115 4.125 78.445 4.295 ;
        RECT 77.960 3.495 78.130 3.955 ;
        RECT 78.430 3.495 78.600 3.955 ;
        RECT 78.115 3.155 78.445 3.325 ;
        RECT 79.000 2.815 79.170 4.635 ;
        RECT 77.390 2.645 79.170 2.815 ;
        RECT 85.200 4.655 86.980 4.825 ;
        RECT 85.200 2.835 85.370 4.655 ;
        RECT 85.925 4.145 86.255 4.315 ;
        RECT 85.770 3.515 85.940 3.975 ;
        RECT 86.240 3.515 86.410 3.975 ;
        RECT 85.925 3.175 86.255 3.345 ;
        RECT 86.810 2.835 86.980 4.655 ;
        RECT 85.200 2.665 86.980 2.835 ;
        RECT 92.790 4.635 94.570 4.805 ;
        RECT 92.790 2.815 92.960 4.635 ;
        RECT 93.515 4.125 93.845 4.295 ;
        RECT 93.360 3.495 93.530 3.955 ;
        RECT 93.830 3.495 94.000 3.955 ;
        RECT 93.515 3.155 93.845 3.325 ;
        RECT 94.400 2.815 94.570 4.635 ;
        RECT 92.790 2.645 94.570 2.815 ;
        RECT 100.180 4.605 101.960 4.775 ;
        RECT 100.180 2.785 100.350 4.605 ;
        RECT 100.905 4.095 101.235 4.265 ;
        RECT 100.750 3.465 100.920 3.925 ;
        RECT 101.220 3.465 101.390 3.925 ;
        RECT 100.905 3.125 101.235 3.295 ;
        RECT 101.790 2.785 101.960 4.605 ;
        RECT 106.640 3.235 106.810 5.055 ;
        RECT 107.365 4.545 107.695 4.715 ;
        RECT 107.210 3.915 107.380 4.375 ;
        RECT 107.680 3.915 107.850 4.375 ;
        RECT 107.365 3.575 107.695 3.745 ;
        RECT 108.250 3.235 108.420 5.055 ;
        RECT 139.045 4.735 139.215 6.145 ;
        RECT 141.615 5.875 141.785 6.145 ;
        RECT 139.555 5.275 139.725 5.605 ;
        RECT 139.895 5.575 140.935 5.745 ;
        RECT 139.895 5.135 140.935 5.305 ;
        RECT 141.105 5.275 141.275 5.605 ;
        RECT 141.615 4.975 141.985 5.875 ;
        RECT 141.615 4.735 141.785 4.975 ;
        RECT 139.045 4.565 141.785 4.735 ;
        RECT 106.640 3.065 108.420 3.235 ;
        RECT 117.935 4.025 122.265 4.195 ;
        RECT 107.030 2.955 108.040 3.065 ;
        RECT 100.180 2.615 101.960 2.785 ;
        RECT 117.935 2.615 118.105 4.025 ;
        RECT 118.445 3.155 118.615 3.485 ;
        RECT 118.830 3.455 121.370 3.625 ;
        RECT 118.830 3.015 121.370 3.185 ;
        RECT 121.585 3.155 121.755 3.485 ;
        RECT 122.095 2.615 122.265 4.025 ;
        RECT 138.285 3.305 142.615 3.475 ;
        RECT 138.285 2.965 138.455 3.305 ;
        RECT 117.935 2.445 122.265 2.615 ;
        RECT 45.410 1.975 47.190 2.145 ;
        RECT 54.200 2.175 55.980 2.345 ;
        RECT 14.080 0.780 30.820 0.950 ;
        RECT 14.080 -0.660 14.250 0.780 ;
        RECT 14.930 0.210 29.970 0.380 ;
        RECT 14.930 -0.260 29.970 -0.090 ;
        RECT 30.650 -0.660 30.820 0.780 ;
        RECT 54.200 0.355 54.370 2.175 ;
        RECT 54.925 1.665 55.255 1.835 ;
        RECT 54.770 1.035 54.940 1.495 ;
        RECT 55.240 1.035 55.410 1.495 ;
        RECT 54.925 0.695 55.255 0.865 ;
        RECT 54.630 0.355 55.580 0.375 ;
        RECT 55.810 0.355 55.980 2.175 ;
        RECT 54.200 0.185 55.980 0.355 ;
        RECT 61.790 2.225 63.570 2.395 ;
        RECT 61.790 0.405 61.960 2.225 ;
        RECT 62.515 1.715 62.845 1.885 ;
        RECT 62.360 1.085 62.530 1.545 ;
        RECT 62.830 1.085 63.000 1.545 ;
        RECT 62.515 0.745 62.845 0.915 ;
        RECT 62.220 0.405 63.170 0.425 ;
        RECT 63.400 0.405 63.570 2.225 ;
        RECT 61.790 0.235 63.570 0.405 ;
        RECT 69.400 2.245 71.180 2.415 ;
        RECT 69.400 0.425 69.570 2.245 ;
        RECT 70.125 1.735 70.455 1.905 ;
        RECT 69.970 1.105 70.140 1.565 ;
        RECT 70.440 1.105 70.610 1.565 ;
        RECT 70.125 0.765 70.455 0.935 ;
        RECT 69.830 0.425 70.780 0.445 ;
        RECT 71.010 0.425 71.180 2.245 ;
        RECT 69.400 0.255 71.180 0.425 ;
        RECT 77.400 2.205 79.180 2.375 ;
        RECT 77.400 0.385 77.570 2.205 ;
        RECT 78.125 1.695 78.455 1.865 ;
        RECT 77.970 1.065 78.140 1.525 ;
        RECT 78.440 1.065 78.610 1.525 ;
        RECT 78.125 0.725 78.455 0.895 ;
        RECT 77.830 0.385 78.780 0.405 ;
        RECT 79.010 0.385 79.180 2.205 ;
        RECT 77.400 0.215 79.180 0.385 ;
        RECT 85.210 2.225 86.990 2.395 ;
        RECT 85.210 0.405 85.380 2.225 ;
        RECT 85.935 1.715 86.265 1.885 ;
        RECT 85.780 1.085 85.950 1.545 ;
        RECT 86.250 1.085 86.420 1.545 ;
        RECT 85.935 0.745 86.265 0.915 ;
        RECT 85.640 0.405 86.590 0.425 ;
        RECT 86.820 0.405 86.990 2.225 ;
        RECT 85.210 0.235 86.990 0.405 ;
        RECT 92.800 2.205 94.580 2.375 ;
        RECT 92.800 0.385 92.970 2.205 ;
        RECT 93.525 1.695 93.855 1.865 ;
        RECT 93.370 1.065 93.540 1.525 ;
        RECT 93.840 1.065 94.010 1.525 ;
        RECT 93.525 0.725 93.855 0.895 ;
        RECT 93.230 0.385 94.180 0.405 ;
        RECT 94.410 0.385 94.580 2.205 ;
        RECT 92.800 0.215 94.580 0.385 ;
        RECT 100.190 2.175 101.970 2.345 ;
        RECT 138.145 2.215 138.455 2.965 ;
        RECT 138.795 2.435 138.965 2.765 ;
        RECT 139.180 2.735 141.720 2.905 ;
        RECT 139.180 2.295 141.720 2.465 ;
        RECT 141.935 2.435 142.105 2.765 ;
        RECT 100.190 0.355 100.360 2.175 ;
        RECT 100.915 1.665 101.245 1.835 ;
        RECT 100.760 1.035 100.930 1.495 ;
        RECT 101.230 1.035 101.400 1.495 ;
        RECT 100.915 0.695 101.245 0.865 ;
        RECT 100.620 0.355 101.570 0.375 ;
        RECT 101.800 0.355 101.970 2.175 ;
        RECT 138.285 1.895 138.455 2.215 ;
        RECT 142.445 1.895 142.615 3.305 ;
        RECT 138.285 1.725 142.615 1.895 ;
        RECT 100.190 0.185 101.970 0.355 ;
        RECT 14.080 -0.830 30.820 -0.660 ;
      LAYER met1 ;
        RECT 68.640 87.180 73.450 87.700 ;
        RECT 68.640 72.900 69.160 87.180 ;
        RECT 68.610 71.900 73.350 72.900 ;
        RECT 68.640 66.760 69.160 71.900 ;
        RECT 77.810 71.870 78.810 72.930 ;
        RECT 68.610 66.240 69.190 66.760 ;
        RECT 61.550 63.910 62.070 63.940 ;
        RECT 61.550 63.390 72.770 63.910 ;
        RECT 61.550 63.360 62.070 63.390 ;
        RECT 68.640 47.480 69.160 62.450 ;
        RECT 64.260 46.960 69.160 47.480 ;
        RECT 72.250 45.450 72.770 63.390 ;
        RECT 57.560 44.930 72.770 45.450 ;
        RECT 57.560 43.730 58.080 44.930 ;
        RECT 57.600 42.830 57.920 43.730 ;
        RECT 57.570 40.725 57.950 42.830 ;
        RECT -5.180 31.900 -4.900 33.280 ;
        RECT -4.610 32.750 13.460 32.980 ;
        RECT 12.110 32.100 12.370 32.750 ;
        RECT 13.870 31.900 14.030 31.920 ;
        RECT 40.480 31.900 40.760 33.250 ;
        RECT -5.180 31.620 40.760 31.900 ;
        RECT 12.080 31.050 13.670 31.310 ;
        RECT 13.870 29.590 14.030 31.620 ;
        RECT 14.660 31.310 14.920 31.340 ;
        RECT 14.660 31.050 25.920 31.310 ;
        RECT 14.660 31.020 14.920 31.050 ;
        RECT 13.790 29.330 14.110 29.590 ;
        RECT 13.820 27.720 14.080 28.040 ;
        RECT 23.695 27.970 23.925 31.050 ;
        RECT 25.740 28.550 25.920 31.050 ;
        RECT 25.740 28.370 26.610 28.550 ;
        RECT 25.740 28.180 25.920 28.370 ;
        RECT 2.470 26.960 2.700 27.135 ;
        RECT 10.130 27.000 10.360 27.185 ;
        RECT 2.470 26.740 3.740 26.960 ;
        RECT 2.470 26.595 2.700 26.740 ;
        RECT 1.100 25.500 1.420 25.520 ;
        RECT 3.520 25.500 3.740 26.740 ;
        RECT 9.090 26.840 10.360 27.000 ;
        RECT 9.090 25.590 9.250 26.840 ;
        RECT 10.130 26.645 10.360 26.840 ;
        RECT 10.600 27.060 10.830 27.185 ;
        RECT 10.600 26.850 11.990 27.060 ;
        RECT 10.600 26.645 10.830 26.850 ;
        RECT 9.700 25.830 11.260 25.930 ;
        RECT 9.500 25.640 11.390 25.830 ;
        RECT 9.500 25.590 11.540 25.640 ;
        RECT 1.100 25.280 6.840 25.500 ;
        RECT 9.090 25.430 11.540 25.590 ;
        RECT 11.220 25.380 11.540 25.430 ;
        RECT 1.100 25.260 1.420 25.280 ;
        RECT 6.620 24.480 6.840 25.280 ;
        RECT 11.780 24.525 11.990 26.850 ;
        RECT 12.440 25.350 12.700 25.670 ;
        RECT 8.355 24.480 11.990 24.525 ;
        RECT 6.620 24.315 11.990 24.480 ;
        RECT 12.490 24.680 12.650 25.350 ;
        RECT 13.870 24.680 14.030 27.720 ;
        RECT 23.680 27.650 23.940 27.970 ;
        RECT 25.700 27.860 25.960 28.180 ;
        RECT 26.430 28.010 26.610 28.370 ;
        RECT 26.300 28.000 27.220 28.010 ;
        RECT 26.300 27.800 27.280 28.000 ;
        RECT 26.585 27.770 27.280 27.800 ;
        RECT 20.640 27.150 22.540 27.400 ;
        RECT 20.645 27.140 20.935 27.150 ;
        RECT 20.440 26.720 20.670 26.935 ;
        RECT 12.490 24.520 14.030 24.680 ;
        RECT 19.340 26.520 20.670 26.720 ;
        RECT 6.620 24.260 8.565 24.315 ;
        RECT 1.100 24.110 1.420 24.130 ;
        RECT 2.020 24.110 2.250 24.240 ;
        RECT 1.100 23.890 2.250 24.110 ;
        RECT 1.100 23.870 1.420 23.890 ;
        RECT 2.020 23.820 2.250 23.890 ;
        RECT 2.490 24.210 2.720 24.240 ;
        RECT 2.490 23.960 3.770 24.210 ;
        RECT 2.490 23.820 2.720 23.960 ;
        RECT 3.520 23.195 3.770 23.960 ;
        RECT 2.605 23.150 3.770 23.195 ;
        RECT 1.510 22.945 3.770 23.150 ;
        RECT 1.510 22.480 3.370 22.945 ;
        RECT 2.240 16.750 2.520 22.480 ;
        RECT 7.700 22.000 7.980 22.030 ;
        RECT 6.850 21.720 7.980 22.000 ;
        RECT 6.850 21.020 7.130 21.720 ;
        RECT 7.700 21.690 7.980 21.720 ;
        RECT 8.355 21.445 8.565 24.260 ;
        RECT 8.790 21.720 10.680 22.000 ;
        RECT 10.150 21.445 10.380 21.580 ;
        RECT 8.355 21.235 10.380 21.445 ;
        RECT 10.150 21.160 10.380 21.235 ;
        RECT 10.620 21.390 10.850 21.580 ;
        RECT 12.490 21.390 12.650 24.520 ;
        RECT 19.340 23.970 19.540 26.520 ;
        RECT 20.440 26.395 20.670 26.520 ;
        RECT 22.290 26.825 22.540 27.150 ;
        RECT 24.550 27.270 26.670 27.510 ;
        RECT 24.550 26.825 24.790 27.270 ;
        RECT 26.355 27.260 26.645 27.270 ;
        RECT 22.290 26.575 24.790 26.825 ;
        RECT 25.670 26.850 25.990 26.890 ;
        RECT 26.150 26.850 26.380 27.055 ;
        RECT 25.670 26.670 26.380 26.850 ;
        RECT 25.670 26.630 25.990 26.670 ;
        RECT 22.290 26.280 22.540 26.575 ;
        RECT 24.550 26.320 24.790 26.575 ;
        RECT 26.150 26.515 26.380 26.670 ;
        RECT 24.550 26.310 26.640 26.320 ;
        RECT 22.290 26.245 22.570 26.280 ;
        RECT 20.655 26.190 22.570 26.245 ;
        RECT 20.645 25.995 22.570 26.190 ;
        RECT 24.550 26.080 26.645 26.310 ;
        RECT 20.645 25.960 20.935 25.995 ;
        RECT 22.370 23.970 22.570 25.995 ;
        RECT 23.680 25.740 23.940 26.060 ;
        RECT 10.620 21.230 12.650 21.390 ;
        RECT 14.920 23.770 22.570 23.970 ;
        RECT 10.620 21.160 10.850 21.230 ;
        RECT 6.850 20.740 10.690 21.020 ;
        RECT 6.850 16.750 7.130 20.740 ;
        RECT 9.720 20.470 11.280 20.490 ;
        RECT 11.790 20.470 11.950 21.230 ;
        RECT 9.720 20.310 11.950 20.470 ;
        RECT 9.720 20.260 11.280 20.310 ;
        RECT 14.920 19.070 15.120 23.770 ;
        RECT 18.260 19.460 18.490 19.565 ;
        RECT 18.730 19.460 18.960 19.565 ;
        RECT 19.300 19.460 19.530 20.370 ;
        RECT 23.695 19.460 23.925 25.740 ;
        RECT 78.090 22.260 78.530 71.870 ;
        RECT 88.510 49.700 137.625 49.970 ;
        RECT 88.510 37.410 88.780 49.700 ;
        RECT 99.985 48.115 103.485 48.185 ;
        RECT 99.985 47.915 130.055 48.115 ;
        RECT 99.985 41.385 100.255 47.915 ;
        RECT 103.110 47.845 130.055 47.915 ;
        RECT 102.975 43.840 103.285 44.270 ;
        RECT 104.650 43.840 104.910 43.900 ;
        RECT 101.525 43.640 104.910 43.840 ;
        RECT 123.075 43.790 124.075 44.820 ;
        RECT 101.525 42.010 101.725 43.640 ;
        RECT 102.975 43.630 103.285 43.640 ;
        RECT 104.650 43.580 104.910 43.640 ;
        RECT 123.365 43.365 123.685 43.790 ;
        RECT 103.735 43.090 107.055 43.290 ;
        RECT 103.735 42.200 103.935 43.090 ;
        RECT 105.205 42.400 105.795 42.710 ;
        RECT 101.525 41.720 101.755 42.010 ;
        RECT 101.960 41.970 104.460 42.200 ;
        RECT 104.650 42.100 104.910 42.400 ;
        RECT 101.525 41.710 101.725 41.720 ;
        RECT 101.960 41.530 104.460 41.760 ;
        RECT 104.615 41.670 104.945 42.100 ;
        RECT 90.935 41.115 100.255 41.385 ;
        RECT 88.050 36.410 89.050 37.410 ;
        RECT 88.470 36.020 88.770 36.410 ;
        RECT 88.040 34.670 89.040 36.020 ;
        RECT 87.040 34.485 87.360 34.500 ;
        RECT 87.640 34.485 89.450 34.670 ;
        RECT 87.040 34.255 89.450 34.485 ;
        RECT 87.040 34.240 87.360 34.255 ;
        RECT 87.640 33.800 89.450 34.255 ;
        RECT 88.440 33.490 88.730 33.500 ;
        RECT 86.450 33.230 88.780 33.490 ;
        RECT 82.360 29.600 83.360 30.600 ;
        RECT 85.140 30.300 86.140 30.600 ;
        RECT 84.720 30.130 86.140 30.300 ;
        RECT 86.450 30.340 86.710 33.230 ;
        RECT 87.040 32.940 87.360 32.955 ;
        RECT 88.250 32.940 88.480 33.065 ;
        RECT 87.040 32.710 88.480 32.940 ;
        RECT 87.040 32.695 87.360 32.710 ;
        RECT 88.250 30.565 88.480 32.710 ;
        RECT 88.690 31.810 88.920 33.065 ;
        RECT 88.690 31.600 90.200 31.810 ;
        RECT 88.690 30.565 88.920 31.600 ;
        RECT 88.440 30.340 88.730 30.360 ;
        RECT 86.450 30.130 88.780 30.340 ;
        RECT 84.720 30.080 88.780 30.130 ;
        RECT 84.720 30.060 86.730 30.080 ;
        RECT 85.140 29.840 86.730 30.060 ;
        RECT 82.680 28.870 82.880 29.600 ;
        RECT 85.140 29.570 86.140 29.840 ;
        RECT 86.450 28.320 86.710 29.840 ;
        RECT 89.945 29.710 90.155 31.600 ;
        RECT 89.940 29.420 90.725 29.710 ;
        RECT 90.935 29.455 91.205 41.115 ;
        RECT 103.055 40.430 103.235 41.530 ;
        RECT 105.205 41.400 106.685 42.400 ;
        RECT 106.855 41.980 107.055 43.090 ;
        RECT 121.780 43.075 125.275 43.365 ;
        RECT 106.840 41.720 109.770 41.980 ;
        RECT 105.205 41.260 105.795 41.400 ;
        RECT 106.855 40.670 107.055 41.720 ;
        RECT 105.105 40.660 107.055 40.670 ;
        RECT 99.000 40.250 103.235 40.430 ;
        RECT 104.895 40.470 107.055 40.660 ;
        RECT 104.895 40.320 105.165 40.470 ;
        RECT 93.315 33.460 94.315 34.490 ;
        RECT 93.645 32.840 93.895 33.460 ;
        RECT 95.325 32.840 95.585 32.860 ;
        RECT 92.115 32.540 95.595 32.840 ;
        RECT 92.155 31.100 92.415 32.540 ;
        RECT 94.585 31.440 94.845 31.760 ;
        RECT 94.615 31.290 94.815 31.440 ;
        RECT 92.155 30.810 92.445 31.100 ;
        RECT 92.650 31.060 95.150 31.290 ;
        RECT 92.155 30.750 92.415 30.810 ;
        RECT 92.650 30.620 95.150 30.850 ;
        RECT 95.325 30.770 95.585 32.540 ;
        RECT 95.935 32.290 96.195 32.350 ;
        RECT 95.935 32.090 97.775 32.290 ;
        RECT 95.935 32.030 96.195 32.090 ;
        RECT 95.850 31.490 96.370 31.660 ;
        RECT 93.725 29.465 93.915 30.620 ;
        RECT 95.850 30.470 97.160 31.490 ;
        RECT 95.850 30.090 96.370 30.470 ;
        RECT 91.470 29.455 93.920 29.465 ;
        RECT 87.470 29.205 87.790 29.230 ;
        RECT 89.945 29.205 90.155 29.420 ;
        RECT 87.470 28.995 90.155 29.205 ;
        RECT 90.935 29.200 93.920 29.455 ;
        RECT 97.575 29.430 97.775 32.090 ;
        RECT 99.000 29.430 99.180 40.250 ;
        RECT 101.315 39.580 102.055 39.830 ;
        RECT 100.525 38.580 102.055 39.580 ;
        RECT 103.055 39.360 103.235 40.250 ;
        RECT 101.315 38.240 102.055 38.580 ;
        RECT 102.315 39.170 102.555 39.180 ;
        RECT 102.315 38.880 102.585 39.170 ;
        RECT 102.745 39.130 103.745 39.360 ;
        RECT 102.315 37.780 102.555 38.880 ;
        RECT 102.745 38.690 103.745 38.920 ;
        RECT 103.885 38.720 104.145 39.220 ;
        RECT 103.155 38.500 103.355 38.690 ;
        RECT 104.915 38.500 105.115 40.320 ;
        RECT 103.155 38.300 105.115 38.500 ;
        RECT 103.855 37.780 104.175 37.790 ;
        RECT 102.315 37.540 104.175 37.780 ;
        RECT 102.595 36.210 103.595 37.540 ;
        RECT 103.855 37.530 104.175 37.540 ;
        RECT 101.615 34.480 102.615 35.520 ;
        RECT 107.015 34.480 108.015 35.710 ;
        RECT 100.765 34.215 101.085 34.240 ;
        RECT 101.335 34.215 103.075 34.480 ;
        RECT 106.715 34.280 108.445 34.480 ;
        RECT 100.765 34.005 103.075 34.215 ;
        RECT 106.445 34.020 108.445 34.280 ;
        RECT 100.765 33.980 101.085 34.005 ;
        RECT 101.335 33.540 103.075 34.005 ;
        RECT 106.715 33.620 108.445 34.020 ;
        RECT 101.945 33.280 102.235 33.300 ;
        RECT 100.265 33.040 102.235 33.280 ;
        RECT 105.510 33.060 107.770 33.360 ;
        RECT 100.265 30.170 100.545 33.040 ;
        RECT 100.765 32.680 101.085 32.705 ;
        RECT 101.755 32.680 101.985 32.865 ;
        RECT 100.765 32.470 101.985 32.680 ;
        RECT 100.765 32.445 101.085 32.470 ;
        RECT 101.755 30.365 101.985 32.470 ;
        RECT 102.195 31.480 102.425 32.865 ;
        RECT 102.195 31.320 103.425 31.480 ;
        RECT 102.195 30.365 102.425 31.320 ;
        RECT 100.265 29.930 102.285 30.170 ;
        RECT 100.265 29.430 100.545 29.930 ;
        RECT 103.265 29.610 103.425 31.320 ;
        RECT 105.510 30.180 105.810 33.060 ;
        RECT 107.205 32.590 107.435 32.855 ;
        RECT 105.975 32.570 106.295 32.580 ;
        RECT 106.485 32.570 107.435 32.590 ;
        RECT 105.975 32.350 107.435 32.570 ;
        RECT 105.975 32.330 106.735 32.350 ;
        RECT 105.975 32.320 106.295 32.330 ;
        RECT 107.205 30.355 107.435 32.350 ;
        RECT 107.645 31.360 107.875 32.855 ;
        RECT 107.645 31.150 109.090 31.360 ;
        RECT 107.645 30.355 107.875 31.150 ;
        RECT 105.510 29.880 107.730 30.180 ;
        RECT 105.510 29.700 105.810 29.880 ;
        RECT 105.390 29.670 105.810 29.700 ;
        RECT 104.090 29.610 105.810 29.670 ;
        RECT 90.935 29.185 91.645 29.200 ;
        RECT 87.470 28.970 87.790 28.995 ;
        RECT 92.010 28.690 92.660 28.990 ;
        RECT 86.450 28.060 88.790 28.320 ;
        RECT 86.470 26.730 86.730 28.060 ;
        RECT 88.420 28.050 88.710 28.060 ;
        RECT 87.470 27.475 87.790 27.500 ;
        RECT 88.230 27.475 88.460 27.890 ;
        RECT 87.470 27.265 88.460 27.475 ;
        RECT 87.470 27.240 87.790 27.265 ;
        RECT 88.230 26.890 88.460 27.265 ;
        RECT 88.670 27.480 88.900 27.890 ;
        RECT 91.180 27.690 92.660 28.690 ;
        RECT 93.725 28.430 93.915 29.200 ;
        RECT 97.560 29.190 100.545 29.430 ;
        RECT 103.255 29.420 105.810 29.610 ;
        RECT 103.255 29.370 104.605 29.420 ;
        RECT 95.785 28.990 97.775 29.190 ;
        RECT 99.000 29.180 99.180 29.190 ;
        RECT 88.670 27.260 89.660 27.480 ;
        RECT 88.670 26.890 88.900 27.260 ;
        RECT 86.470 26.470 88.730 26.730 ;
        RECT 89.430 26.220 89.650 27.260 ;
        RECT 92.010 27.220 92.660 27.690 ;
        RECT 92.950 28.240 93.140 28.265 ;
        RECT 92.950 27.950 93.185 28.240 ;
        RECT 93.345 28.200 94.345 28.430 ;
        RECT 92.950 26.795 93.140 27.950 ;
        RECT 93.345 27.760 94.345 27.990 ;
        RECT 94.505 27.970 94.735 28.240 ;
        RECT 93.775 27.390 93.975 27.760 ;
        RECT 94.490 27.650 94.750 27.970 ;
        RECT 95.785 27.730 95.985 28.990 ;
        RECT 100.265 28.550 100.545 29.190 ;
        RECT 101.225 29.220 101.545 29.270 ;
        RECT 103.265 29.220 103.425 29.370 ;
        RECT 101.225 29.060 103.425 29.220 ;
        RECT 104.090 29.190 104.605 29.370 ;
        RECT 101.225 29.010 101.545 29.060 ;
        RECT 100.265 28.310 102.295 28.550 ;
        RECT 100.285 28.270 102.295 28.310 ;
        RECT 95.785 27.640 95.995 27.730 ;
        RECT 95.795 27.390 95.995 27.640 ;
        RECT 93.775 27.190 95.995 27.390 ;
        RECT 100.295 26.950 100.585 28.270 ;
        RECT 101.975 28.260 102.265 28.270 ;
        RECT 101.225 27.760 101.545 27.810 ;
        RECT 101.785 27.760 102.015 28.100 ;
        RECT 101.225 27.600 102.015 27.760 ;
        RECT 101.225 27.550 101.545 27.600 ;
        RECT 101.785 27.100 102.015 27.600 ;
        RECT 102.225 27.710 102.455 28.100 ;
        RECT 102.225 27.510 103.115 27.710 ;
        RECT 102.225 27.100 102.455 27.510 ;
        RECT 94.490 26.795 94.750 26.860 ;
        RECT 92.950 26.605 94.750 26.795 ;
        RECT 100.295 26.670 102.315 26.950 ;
        RECT 87.660 25.900 89.650 26.220 ;
        RECT 93.745 25.980 93.965 26.605 ;
        RECT 94.490 26.540 94.750 26.605 ;
        RECT 102.855 26.420 103.055 27.510 ;
        RECT 101.285 26.220 103.055 26.420 ;
        RECT 87.660 25.640 89.440 25.900 ;
        RECT 101.285 25.760 103.045 26.220 ;
        RECT 88.040 24.650 89.040 25.640 ;
        RECT 101.615 25.020 102.615 25.760 ;
        RECT 88.400 24.320 88.680 24.650 ;
        RECT 88.020 23.320 89.020 24.320 ;
        RECT 104.355 24.095 104.605 29.190 ;
        RECT 105.510 28.170 105.810 29.420 ;
        RECT 108.875 29.460 109.085 31.150 ;
        RECT 109.510 29.460 109.770 41.720 ;
        RECT 121.780 41.290 122.070 43.075 ;
        RECT 124.205 42.320 127.805 42.540 ;
        RECT 124.205 41.480 124.425 42.320 ;
        RECT 125.605 41.690 126.405 42.110 ;
        RECT 121.780 41.000 122.105 41.290 ;
        RECT 122.310 41.250 124.810 41.480 ;
        RECT 121.780 40.955 122.070 41.000 ;
        RECT 122.310 40.810 124.810 41.040 ;
        RECT 124.955 40.970 125.245 41.650 ;
        RECT 123.345 39.840 123.545 40.810 ;
        RECT 125.605 40.690 127.265 41.690 ;
        RECT 127.585 41.495 127.805 42.320 ;
        RECT 127.585 41.225 129.355 41.495 ;
        RECT 125.605 40.410 126.405 40.690 ;
        RECT 118.190 39.640 123.545 39.840 ;
        RECT 127.585 39.790 127.805 41.225 ;
        RECT 113.305 33.420 113.615 34.060 ;
        RECT 111.905 33.120 115.355 33.420 ;
        RECT 111.905 31.260 112.205 33.120 ;
        RECT 114.605 32.610 117.375 32.790 ;
        RECT 114.605 31.770 114.785 32.610 ;
        RECT 115.595 32.020 116.455 32.300 ;
        RECT 112.350 31.540 114.850 31.770 ;
        RECT 112.350 31.100 114.850 31.330 ;
        RECT 115.025 31.290 115.325 31.850 ;
        RECT 113.255 30.005 113.435 31.100 ;
        RECT 115.595 31.020 117.035 32.020 ;
        RECT 115.595 30.590 116.455 31.020 ;
        RECT 117.195 30.420 117.375 32.610 ;
        RECT 118.190 30.420 118.390 39.640 ;
        RECT 121.915 38.820 122.325 39.160 ;
        RECT 120.985 37.820 122.325 38.820 ;
        RECT 123.345 38.610 123.545 39.640 ;
        RECT 125.195 39.570 127.805 39.790 ;
        RECT 122.565 38.420 122.770 38.470 ;
        RECT 122.545 38.130 122.775 38.420 ;
        RECT 122.935 38.380 123.935 38.610 ;
        RECT 121.915 37.400 122.325 37.820 ;
        RECT 122.565 37.110 122.770 38.130 ;
        RECT 122.935 37.940 123.935 38.170 ;
        RECT 123.385 37.660 123.605 37.940 ;
        RECT 124.085 37.830 124.365 38.440 ;
        RECT 125.195 37.660 125.415 39.570 ;
        RECT 123.385 37.440 125.415 37.660 ;
        RECT 122.525 36.830 124.395 37.110 ;
        RECT 123.205 36.190 123.555 36.830 ;
        RECT 119.350 34.590 119.670 34.625 ;
        RECT 120.315 34.620 121.315 36.180 ;
        RECT 119.955 34.590 121.775 34.620 ;
        RECT 119.350 34.400 121.775 34.590 ;
        RECT 125.385 34.570 126.385 35.960 ;
        RECT 125.025 34.560 126.865 34.570 ;
        RECT 119.350 34.365 119.670 34.400 ;
        RECT 119.955 33.930 121.775 34.400 ;
        RECT 124.225 34.300 126.865 34.560 ;
        RECT 125.025 33.710 126.865 34.300 ;
        RECT 118.970 33.380 121.050 33.660 ;
        RECT 118.970 32.710 119.250 33.380 ;
        RECT 123.605 33.270 126.125 33.570 ;
        RECT 118.970 32.080 119.210 32.710 ;
        RECT 119.380 32.475 119.640 32.540 ;
        RECT 120.565 32.475 120.795 33.225 ;
        RECT 119.380 32.285 120.795 32.475 ;
        RECT 119.380 32.220 119.640 32.285 ;
        RECT 118.970 30.500 119.250 32.080 ;
        RECT 120.565 30.725 120.795 32.285 ;
        RECT 121.005 32.020 121.235 33.225 ;
        RECT 123.605 32.130 123.905 33.270 ;
        RECT 125.775 33.200 126.065 33.270 ;
        RECT 125.585 32.610 125.815 32.995 ;
        RECT 124.225 32.350 125.815 32.610 ;
        RECT 121.005 31.770 122.315 32.020 ;
        RECT 123.605 31.830 124.635 32.130 ;
        RECT 121.005 30.725 121.235 31.770 ;
        RECT 120.755 30.500 121.045 30.520 ;
        RECT 118.970 30.420 121.120 30.500 ;
        RECT 117.185 30.240 121.120 30.420 ;
        RECT 115.415 30.220 121.120 30.240 ;
        RECT 115.415 30.190 119.320 30.220 ;
        RECT 115.415 30.060 117.375 30.190 ;
        RECT 108.875 29.200 109.770 29.460 ;
        RECT 110.615 29.755 113.465 30.005 ;
        RECT 106.690 29.075 107.010 29.100 ;
        RECT 108.875 29.075 109.085 29.200 ;
        RECT 106.690 28.865 109.085 29.075 ;
        RECT 106.690 28.840 107.010 28.865 ;
        RECT 105.510 27.870 107.830 28.170 ;
        RECT 105.510 26.560 105.810 27.870 ;
        RECT 106.690 27.395 107.010 27.420 ;
        RECT 107.265 27.395 107.495 27.720 ;
        RECT 106.690 27.185 107.495 27.395 ;
        RECT 106.690 27.160 107.010 27.185 ;
        RECT 107.265 26.720 107.495 27.185 ;
        RECT 107.705 27.350 107.935 27.720 ;
        RECT 107.705 27.110 108.615 27.350 ;
        RECT 107.705 26.720 107.935 27.110 ;
        RECT 105.510 26.260 107.820 26.560 ;
        RECT 108.375 26.020 108.615 27.110 ;
        RECT 106.640 25.690 108.615 26.020 ;
        RECT 106.640 25.420 108.530 25.690 ;
        RECT 107.250 24.600 108.250 25.420 ;
        RECT 110.615 24.095 110.865 29.755 ;
        RECT 111.885 29.130 112.475 29.580 ;
        RECT 111.145 28.130 112.475 29.130 ;
        RECT 113.255 29.010 113.435 29.755 ;
        RECT 111.885 27.780 112.475 28.130 ;
        RECT 112.735 27.490 112.985 28.850 ;
        RECT 113.145 28.780 114.145 29.010 ;
        RECT 114.315 28.820 114.555 28.830 ;
        RECT 113.145 28.340 114.145 28.570 ;
        RECT 114.305 28.530 114.555 28.820 ;
        RECT 113.535 27.940 113.715 28.340 ;
        RECT 114.305 28.210 114.565 28.530 ;
        RECT 114.315 28.180 114.555 28.210 ;
        RECT 115.415 27.940 115.595 30.060 ;
        RECT 113.535 27.760 115.595 27.940 ;
        RECT 118.970 28.840 119.250 30.190 ;
        RECT 122.060 30.140 122.310 31.770 ;
        RECT 124.335 30.320 124.635 31.830 ;
        RECT 125.585 30.495 125.815 32.350 ;
        RECT 126.025 31.730 126.255 32.995 ;
        RECT 126.025 31.470 127.525 31.730 ;
        RECT 126.025 30.495 126.255 31.470 ;
        RECT 124.325 30.210 126.145 30.320 ;
        RECT 123.585 30.140 126.145 30.210 ;
        RECT 122.060 30.020 126.145 30.140 ;
        RECT 122.060 29.940 124.635 30.020 ;
        RECT 122.060 29.910 123.835 29.940 ;
        RECT 119.755 29.655 120.075 29.660 ;
        RECT 122.060 29.655 122.310 29.910 ;
        RECT 119.755 29.405 122.310 29.655 ;
        RECT 119.755 29.400 120.075 29.405 ;
        RECT 118.970 28.560 121.100 28.840 ;
        RECT 112.725 27.230 112.985 27.490 ;
        RECT 114.275 27.300 114.595 27.560 ;
        RECT 112.725 27.080 112.965 27.230 ;
        RECT 114.315 27.080 114.555 27.300 ;
        RECT 112.725 26.840 114.555 27.080 ;
        RECT 118.970 27.180 119.250 28.560 ;
        RECT 120.785 28.520 121.075 28.560 ;
        RECT 119.785 27.965 120.045 28.000 ;
        RECT 120.595 27.965 120.825 28.360 ;
        RECT 119.785 27.715 120.825 27.965 ;
        RECT 121.035 27.930 121.265 28.360 ;
        RECT 119.785 27.680 120.045 27.715 ;
        RECT 120.595 27.360 120.825 27.715 ;
        RECT 120.995 27.650 122.105 27.930 ;
        RECT 121.035 27.360 121.265 27.650 ;
        RECT 120.785 27.180 121.075 27.200 ;
        RECT 118.970 26.970 121.075 27.180 ;
        RECT 118.970 26.900 121.060 26.970 ;
        RECT 112.855 26.500 114.405 26.840 ;
        RECT 121.825 26.710 122.105 27.650 ;
        RECT 113.165 25.620 114.165 26.500 ;
        RECT 119.985 26.250 122.105 26.710 ;
        RECT 119.985 25.930 121.825 26.250 ;
        RECT 120.665 25.130 121.665 25.930 ;
        RECT 104.355 23.845 110.865 24.095 ;
        RECT 123.070 24.270 123.290 29.910 ;
        RECT 124.325 28.520 124.625 29.940 ;
        RECT 127.265 29.900 127.525 31.470 ;
        RECT 129.085 29.900 129.355 41.225 ;
        RECT 129.785 29.900 130.055 47.845 ;
        RECT 137.355 44.515 137.625 49.700 ;
        RECT 148.920 47.745 152.420 47.815 ;
        RECT 148.920 47.545 178.990 47.745 ;
        RECT 137.355 44.185 138.705 44.515 ;
        RECT 137.355 35.650 137.625 44.185 ;
        RECT 148.920 41.015 149.190 47.545 ;
        RECT 152.045 47.475 178.990 47.545 ;
        RECT 151.910 43.470 152.220 43.900 ;
        RECT 153.585 43.470 153.845 43.530 ;
        RECT 150.460 43.270 153.845 43.470 ;
        RECT 172.010 43.420 173.010 44.450 ;
        RECT 150.460 41.640 150.660 43.270 ;
        RECT 151.910 43.260 152.220 43.270 ;
        RECT 153.585 43.210 153.845 43.270 ;
        RECT 172.300 42.995 172.620 43.420 ;
        RECT 152.670 42.720 155.990 42.920 ;
        RECT 152.670 41.830 152.870 42.720 ;
        RECT 154.140 42.030 154.730 42.340 ;
        RECT 150.460 41.350 150.690 41.640 ;
        RECT 150.895 41.600 153.395 41.830 ;
        RECT 153.585 41.730 153.845 42.030 ;
        RECT 150.460 41.340 150.660 41.350 ;
        RECT 150.895 41.160 153.395 41.390 ;
        RECT 153.550 41.300 153.880 41.730 ;
        RECT 139.870 40.745 149.190 41.015 ;
        RECT 136.975 34.300 137.975 35.650 ;
        RECT 135.975 34.115 136.295 34.130 ;
        RECT 136.575 34.115 138.385 34.300 ;
        RECT 135.975 33.885 138.385 34.115 ;
        RECT 135.975 33.870 136.295 33.885 ;
        RECT 136.575 33.430 138.385 33.885 ;
        RECT 137.375 33.120 137.665 33.130 ;
        RECT 135.385 32.860 137.715 33.120 ;
        RECT 127.265 29.630 131.725 29.900 ;
        RECT 134.075 29.760 135.075 30.230 ;
        RECT 135.385 29.970 135.645 32.860 ;
        RECT 135.975 32.570 136.295 32.585 ;
        RECT 137.185 32.570 137.415 32.695 ;
        RECT 135.975 32.340 137.415 32.570 ;
        RECT 135.975 32.325 136.295 32.340 ;
        RECT 137.185 30.195 137.415 32.340 ;
        RECT 137.625 31.440 137.855 32.695 ;
        RECT 137.625 31.230 139.135 31.440 ;
        RECT 137.625 30.195 137.855 31.230 ;
        RECT 137.375 29.970 137.665 29.990 ;
        RECT 135.385 29.760 137.715 29.970 ;
        RECT 134.075 29.720 137.715 29.760 ;
        RECT 133.900 29.710 137.715 29.720 ;
        RECT 127.265 29.420 127.525 29.630 ;
        RECT 124.895 29.160 127.525 29.420 ;
        RECT 133.900 29.470 135.665 29.710 ;
        RECT 133.900 29.200 135.075 29.470 ;
        RECT 133.900 28.760 134.120 29.200 ;
        RECT 128.500 28.540 134.120 28.760 ;
        RECT 124.255 28.450 126.085 28.520 ;
        RECT 124.255 28.220 126.095 28.450 ;
        RECT 124.325 26.900 124.625 28.220 ;
        RECT 125.615 27.680 125.845 28.060 ;
        RECT 124.895 27.420 125.845 27.680 ;
        RECT 125.615 27.060 125.845 27.420 ;
        RECT 126.055 27.330 126.285 28.060 ;
        RECT 126.055 27.140 126.955 27.330 ;
        RECT 126.055 27.060 126.285 27.140 ;
        RECT 124.325 26.890 125.405 26.900 ;
        RECT 125.805 26.890 126.095 26.900 ;
        RECT 124.325 26.650 126.155 26.890 ;
        RECT 126.765 26.340 126.955 27.140 ;
        RECT 124.995 26.045 126.955 26.340 ;
        RECT 124.995 25.710 126.895 26.045 ;
        RECT 125.495 24.530 126.495 25.710 ;
        RECT 128.500 24.270 128.720 28.540 ;
        RECT 135.385 27.950 135.645 29.470 ;
        RECT 138.880 29.340 139.090 31.230 ;
        RECT 138.875 29.050 139.660 29.340 ;
        RECT 139.870 29.085 140.140 40.745 ;
        RECT 151.990 40.060 152.170 41.160 ;
        RECT 154.140 41.030 155.620 42.030 ;
        RECT 155.790 41.610 155.990 42.720 ;
        RECT 170.715 42.705 174.210 42.995 ;
        RECT 155.775 41.350 158.705 41.610 ;
        RECT 154.140 40.890 154.730 41.030 ;
        RECT 155.790 40.300 155.990 41.350 ;
        RECT 154.040 40.290 155.990 40.300 ;
        RECT 147.935 39.880 152.170 40.060 ;
        RECT 153.830 40.100 155.990 40.290 ;
        RECT 153.830 39.950 154.100 40.100 ;
        RECT 142.250 33.090 143.250 34.120 ;
        RECT 142.580 32.470 142.830 33.090 ;
        RECT 144.260 32.470 144.520 32.490 ;
        RECT 141.050 32.170 144.530 32.470 ;
        RECT 141.090 30.730 141.350 32.170 ;
        RECT 143.520 31.070 143.780 31.390 ;
        RECT 143.550 30.920 143.750 31.070 ;
        RECT 141.090 30.440 141.380 30.730 ;
        RECT 141.585 30.690 144.085 30.920 ;
        RECT 141.090 30.380 141.350 30.440 ;
        RECT 141.585 30.250 144.085 30.480 ;
        RECT 144.260 30.400 144.520 32.170 ;
        RECT 144.870 31.920 145.130 31.980 ;
        RECT 144.870 31.720 146.710 31.920 ;
        RECT 144.870 31.660 145.130 31.720 ;
        RECT 144.785 31.120 145.305 31.290 ;
        RECT 142.660 29.095 142.850 30.250 ;
        RECT 144.785 30.100 146.095 31.120 ;
        RECT 144.785 29.720 145.305 30.100 ;
        RECT 140.405 29.085 142.855 29.095 ;
        RECT 136.405 28.835 136.725 28.860 ;
        RECT 138.880 28.835 139.090 29.050 ;
        RECT 136.405 28.625 139.090 28.835 ;
        RECT 139.870 28.830 142.855 29.085 ;
        RECT 146.510 29.060 146.710 31.720 ;
        RECT 147.935 29.060 148.115 39.880 ;
        RECT 150.250 39.210 150.990 39.460 ;
        RECT 149.460 38.210 150.990 39.210 ;
        RECT 151.990 38.990 152.170 39.880 ;
        RECT 150.250 37.870 150.990 38.210 ;
        RECT 151.250 38.800 151.490 38.810 ;
        RECT 151.250 38.510 151.520 38.800 ;
        RECT 151.680 38.760 152.680 38.990 ;
        RECT 151.250 37.410 151.490 38.510 ;
        RECT 151.680 38.320 152.680 38.550 ;
        RECT 152.820 38.350 153.080 38.850 ;
        RECT 152.090 38.130 152.290 38.320 ;
        RECT 153.850 38.130 154.050 39.950 ;
        RECT 152.090 37.930 154.050 38.130 ;
        RECT 152.790 37.410 153.110 37.420 ;
        RECT 151.250 37.170 153.110 37.410 ;
        RECT 151.530 35.840 152.530 37.170 ;
        RECT 152.790 37.160 153.110 37.170 ;
        RECT 150.550 34.110 151.550 35.150 ;
        RECT 155.950 34.110 156.950 35.340 ;
        RECT 149.700 33.845 150.020 33.870 ;
        RECT 150.270 33.845 152.010 34.110 ;
        RECT 155.650 33.910 157.380 34.110 ;
        RECT 149.700 33.635 152.010 33.845 ;
        RECT 155.380 33.650 157.380 33.910 ;
        RECT 149.700 33.610 150.020 33.635 ;
        RECT 150.270 33.170 152.010 33.635 ;
        RECT 155.650 33.250 157.380 33.650 ;
        RECT 150.880 32.910 151.170 32.930 ;
        RECT 149.200 32.670 151.170 32.910 ;
        RECT 154.445 32.690 156.705 32.990 ;
        RECT 149.200 29.800 149.480 32.670 ;
        RECT 149.700 32.310 150.020 32.335 ;
        RECT 150.690 32.310 150.920 32.495 ;
        RECT 149.700 32.100 150.920 32.310 ;
        RECT 149.700 32.075 150.020 32.100 ;
        RECT 150.690 29.995 150.920 32.100 ;
        RECT 151.130 31.110 151.360 32.495 ;
        RECT 151.130 30.950 152.360 31.110 ;
        RECT 151.130 29.995 151.360 30.950 ;
        RECT 149.200 29.560 151.220 29.800 ;
        RECT 149.200 29.060 149.480 29.560 ;
        RECT 152.200 29.240 152.360 30.950 ;
        RECT 154.445 29.810 154.745 32.690 ;
        RECT 156.140 32.220 156.370 32.485 ;
        RECT 154.910 32.200 155.230 32.210 ;
        RECT 155.420 32.200 156.370 32.220 ;
        RECT 154.910 31.980 156.370 32.200 ;
        RECT 154.910 31.960 155.670 31.980 ;
        RECT 154.910 31.950 155.230 31.960 ;
        RECT 156.140 29.985 156.370 31.980 ;
        RECT 156.580 30.990 156.810 32.485 ;
        RECT 156.580 30.780 158.025 30.990 ;
        RECT 156.580 29.985 156.810 30.780 ;
        RECT 154.445 29.510 156.665 29.810 ;
        RECT 154.445 29.330 154.745 29.510 ;
        RECT 154.325 29.300 154.745 29.330 ;
        RECT 153.025 29.240 154.745 29.300 ;
        RECT 139.870 28.815 140.580 28.830 ;
        RECT 136.405 28.600 136.725 28.625 ;
        RECT 140.945 28.320 141.595 28.620 ;
        RECT 135.385 27.690 137.725 27.950 ;
        RECT 135.405 26.360 135.665 27.690 ;
        RECT 137.355 27.680 137.645 27.690 ;
        RECT 136.405 27.105 136.725 27.130 ;
        RECT 137.165 27.105 137.395 27.520 ;
        RECT 136.405 26.895 137.395 27.105 ;
        RECT 136.405 26.870 136.725 26.895 ;
        RECT 137.165 26.520 137.395 26.895 ;
        RECT 137.605 27.110 137.835 27.520 ;
        RECT 140.115 27.320 141.595 28.320 ;
        RECT 142.660 28.060 142.850 28.830 ;
        RECT 146.495 28.820 149.480 29.060 ;
        RECT 152.190 29.050 154.745 29.240 ;
        RECT 152.190 29.000 153.540 29.050 ;
        RECT 144.720 28.620 146.710 28.820 ;
        RECT 147.935 28.810 148.115 28.820 ;
        RECT 137.605 26.890 138.595 27.110 ;
        RECT 137.605 26.520 137.835 26.890 ;
        RECT 135.405 26.100 137.665 26.360 ;
        RECT 138.365 25.850 138.585 26.890 ;
        RECT 140.945 26.850 141.595 27.320 ;
        RECT 141.885 27.870 142.075 27.895 ;
        RECT 141.885 27.580 142.120 27.870 ;
        RECT 142.280 27.830 143.280 28.060 ;
        RECT 141.885 26.425 142.075 27.580 ;
        RECT 142.280 27.390 143.280 27.620 ;
        RECT 143.440 27.600 143.670 27.870 ;
        RECT 142.710 27.020 142.910 27.390 ;
        RECT 143.425 27.280 143.685 27.600 ;
        RECT 144.720 27.360 144.920 28.620 ;
        RECT 149.200 28.180 149.480 28.820 ;
        RECT 150.160 28.850 150.480 28.900 ;
        RECT 152.200 28.850 152.360 29.000 ;
        RECT 150.160 28.690 152.360 28.850 ;
        RECT 153.025 28.820 153.540 29.000 ;
        RECT 150.160 28.640 150.480 28.690 ;
        RECT 149.200 27.940 151.230 28.180 ;
        RECT 149.220 27.900 151.230 27.940 ;
        RECT 144.720 27.270 144.930 27.360 ;
        RECT 144.730 27.020 144.930 27.270 ;
        RECT 142.710 26.820 144.930 27.020 ;
        RECT 149.230 26.580 149.520 27.900 ;
        RECT 150.910 27.890 151.200 27.900 ;
        RECT 150.160 27.390 150.480 27.440 ;
        RECT 150.720 27.390 150.950 27.730 ;
        RECT 150.160 27.230 150.950 27.390 ;
        RECT 150.160 27.180 150.480 27.230 ;
        RECT 150.720 26.730 150.950 27.230 ;
        RECT 151.160 27.340 151.390 27.730 ;
        RECT 151.160 27.140 152.050 27.340 ;
        RECT 151.160 26.730 151.390 27.140 ;
        RECT 143.425 26.425 143.685 26.490 ;
        RECT 141.885 26.235 143.685 26.425 ;
        RECT 149.230 26.300 151.250 26.580 ;
        RECT 136.595 25.530 138.585 25.850 ;
        RECT 142.680 25.610 142.900 26.235 ;
        RECT 143.425 26.170 143.685 26.235 ;
        RECT 151.790 26.050 151.990 27.140 ;
        RECT 150.220 25.850 151.990 26.050 ;
        RECT 136.595 25.270 138.375 25.530 ;
        RECT 150.220 25.390 151.980 25.850 ;
        RECT 136.975 24.280 137.975 25.270 ;
        RECT 150.550 24.650 151.550 25.390 ;
        RECT 123.070 24.050 128.720 24.270 ;
        RECT 18.260 19.230 23.925 19.460 ;
        RECT 47.300 21.820 78.530 22.260 ;
        RECT 88.350 22.520 88.670 23.320 ;
        RECT 137.380 22.520 137.700 24.280 ;
        RECT 153.290 23.725 153.540 28.820 ;
        RECT 154.445 27.800 154.745 29.050 ;
        RECT 157.810 29.090 158.020 30.780 ;
        RECT 158.445 29.090 158.705 41.350 ;
        RECT 170.715 40.920 171.005 42.705 ;
        RECT 173.140 41.950 176.740 42.170 ;
        RECT 173.140 41.110 173.360 41.950 ;
        RECT 174.540 41.320 175.340 41.740 ;
        RECT 170.715 40.630 171.040 40.920 ;
        RECT 171.245 40.880 173.745 41.110 ;
        RECT 170.715 40.585 171.005 40.630 ;
        RECT 171.245 40.440 173.745 40.670 ;
        RECT 173.890 40.600 174.180 41.280 ;
        RECT 172.280 39.470 172.480 40.440 ;
        RECT 174.540 40.320 176.200 41.320 ;
        RECT 176.520 41.125 176.740 41.950 ;
        RECT 176.520 40.855 178.290 41.125 ;
        RECT 174.540 40.040 175.340 40.320 ;
        RECT 167.125 39.270 172.480 39.470 ;
        RECT 176.520 39.420 176.740 40.855 ;
        RECT 162.240 33.050 162.550 33.690 ;
        RECT 160.840 32.750 164.290 33.050 ;
        RECT 160.840 30.890 161.140 32.750 ;
        RECT 163.540 32.240 166.310 32.420 ;
        RECT 163.540 31.400 163.720 32.240 ;
        RECT 164.530 31.650 165.390 31.930 ;
        RECT 161.285 31.170 163.785 31.400 ;
        RECT 161.285 30.730 163.785 30.960 ;
        RECT 163.960 30.920 164.260 31.480 ;
        RECT 162.190 29.635 162.370 30.730 ;
        RECT 164.530 30.650 165.970 31.650 ;
        RECT 164.530 30.220 165.390 30.650 ;
        RECT 166.130 30.050 166.310 32.240 ;
        RECT 167.125 30.050 167.325 39.270 ;
        RECT 170.850 38.450 171.260 38.790 ;
        RECT 169.920 37.450 171.260 38.450 ;
        RECT 172.280 38.240 172.480 39.270 ;
        RECT 174.130 39.200 176.740 39.420 ;
        RECT 171.500 38.050 171.705 38.100 ;
        RECT 171.480 37.760 171.710 38.050 ;
        RECT 171.870 38.010 172.870 38.240 ;
        RECT 170.850 37.030 171.260 37.450 ;
        RECT 171.500 36.740 171.705 37.760 ;
        RECT 171.870 37.570 172.870 37.800 ;
        RECT 172.320 37.290 172.540 37.570 ;
        RECT 173.020 37.460 173.300 38.070 ;
        RECT 174.130 37.290 174.350 39.200 ;
        RECT 172.320 37.070 174.350 37.290 ;
        RECT 171.460 36.460 173.330 36.740 ;
        RECT 172.140 35.820 172.490 36.460 ;
        RECT 168.285 34.220 168.605 34.255 ;
        RECT 169.250 34.250 170.250 35.810 ;
        RECT 168.890 34.220 170.710 34.250 ;
        RECT 168.285 34.030 170.710 34.220 ;
        RECT 174.320 34.200 175.320 35.590 ;
        RECT 173.960 34.190 175.800 34.200 ;
        RECT 168.285 33.995 168.605 34.030 ;
        RECT 168.890 33.560 170.710 34.030 ;
        RECT 173.160 33.930 175.800 34.190 ;
        RECT 173.960 33.340 175.800 33.930 ;
        RECT 167.905 33.010 169.985 33.290 ;
        RECT 167.905 32.340 168.185 33.010 ;
        RECT 172.540 32.900 175.060 33.200 ;
        RECT 167.905 31.710 168.145 32.340 ;
        RECT 168.315 32.105 168.575 32.170 ;
        RECT 169.500 32.105 169.730 32.855 ;
        RECT 168.315 31.915 169.730 32.105 ;
        RECT 168.315 31.850 168.575 31.915 ;
        RECT 167.905 30.130 168.185 31.710 ;
        RECT 169.500 30.355 169.730 31.915 ;
        RECT 169.940 31.650 170.170 32.855 ;
        RECT 172.540 31.760 172.840 32.900 ;
        RECT 174.710 32.830 175.000 32.900 ;
        RECT 174.520 32.240 174.750 32.625 ;
        RECT 173.160 31.980 174.750 32.240 ;
        RECT 169.940 31.400 171.250 31.650 ;
        RECT 172.540 31.460 173.570 31.760 ;
        RECT 169.940 30.355 170.170 31.400 ;
        RECT 169.690 30.130 169.980 30.150 ;
        RECT 167.905 30.050 170.055 30.130 ;
        RECT 166.120 29.870 170.055 30.050 ;
        RECT 164.350 29.850 170.055 29.870 ;
        RECT 164.350 29.820 168.255 29.850 ;
        RECT 164.350 29.690 166.310 29.820 ;
        RECT 157.810 28.830 158.705 29.090 ;
        RECT 159.550 29.385 162.400 29.635 ;
        RECT 155.625 28.705 155.945 28.730 ;
        RECT 157.810 28.705 158.020 28.830 ;
        RECT 155.625 28.495 158.020 28.705 ;
        RECT 155.625 28.470 155.945 28.495 ;
        RECT 154.445 27.500 156.765 27.800 ;
        RECT 154.445 26.190 154.745 27.500 ;
        RECT 155.625 27.025 155.945 27.050 ;
        RECT 156.200 27.025 156.430 27.350 ;
        RECT 155.625 26.815 156.430 27.025 ;
        RECT 155.625 26.790 155.945 26.815 ;
        RECT 156.200 26.350 156.430 26.815 ;
        RECT 156.640 26.980 156.870 27.350 ;
        RECT 156.640 26.740 157.550 26.980 ;
        RECT 156.640 26.350 156.870 26.740 ;
        RECT 154.445 25.890 156.755 26.190 ;
        RECT 157.310 25.650 157.550 26.740 ;
        RECT 155.575 25.320 157.550 25.650 ;
        RECT 155.575 25.050 157.465 25.320 ;
        RECT 156.185 24.230 157.185 25.050 ;
        RECT 159.550 23.725 159.800 29.385 ;
        RECT 160.820 28.760 161.410 29.210 ;
        RECT 160.080 27.760 161.410 28.760 ;
        RECT 162.190 28.640 162.370 29.385 ;
        RECT 160.820 27.410 161.410 27.760 ;
        RECT 161.670 27.120 161.920 28.480 ;
        RECT 162.080 28.410 163.080 28.640 ;
        RECT 163.250 28.450 163.490 28.460 ;
        RECT 162.080 27.970 163.080 28.200 ;
        RECT 163.240 28.160 163.490 28.450 ;
        RECT 162.470 27.570 162.650 27.970 ;
        RECT 163.240 27.840 163.500 28.160 ;
        RECT 163.250 27.810 163.490 27.840 ;
        RECT 164.350 27.570 164.530 29.690 ;
        RECT 162.470 27.390 164.530 27.570 ;
        RECT 167.905 28.470 168.185 29.820 ;
        RECT 170.995 29.770 171.245 31.400 ;
        RECT 173.270 29.950 173.570 31.460 ;
        RECT 174.520 30.125 174.750 31.980 ;
        RECT 174.960 31.360 175.190 32.625 ;
        RECT 174.960 31.100 176.460 31.360 ;
        RECT 174.960 30.125 175.190 31.100 ;
        RECT 173.260 29.840 175.080 29.950 ;
        RECT 172.520 29.770 175.080 29.840 ;
        RECT 170.995 29.650 175.080 29.770 ;
        RECT 170.995 29.570 173.570 29.650 ;
        RECT 170.995 29.540 172.770 29.570 ;
        RECT 168.690 29.285 169.010 29.290 ;
        RECT 170.995 29.285 171.245 29.540 ;
        RECT 168.690 29.035 171.245 29.285 ;
        RECT 168.690 29.030 169.010 29.035 ;
        RECT 167.905 28.190 170.035 28.470 ;
        RECT 161.660 26.860 161.920 27.120 ;
        RECT 163.210 26.930 163.530 27.190 ;
        RECT 161.660 26.710 161.900 26.860 ;
        RECT 163.250 26.710 163.490 26.930 ;
        RECT 161.660 26.470 163.490 26.710 ;
        RECT 167.905 26.810 168.185 28.190 ;
        RECT 169.720 28.150 170.010 28.190 ;
        RECT 168.720 27.595 168.980 27.630 ;
        RECT 169.530 27.595 169.760 27.990 ;
        RECT 168.720 27.345 169.760 27.595 ;
        RECT 169.970 27.560 170.200 27.990 ;
        RECT 168.720 27.310 168.980 27.345 ;
        RECT 169.530 26.990 169.760 27.345 ;
        RECT 169.930 27.280 171.040 27.560 ;
        RECT 169.970 26.990 170.200 27.280 ;
        RECT 169.720 26.810 170.010 26.830 ;
        RECT 167.905 26.600 170.010 26.810 ;
        RECT 167.905 26.530 169.995 26.600 ;
        RECT 161.790 26.130 163.340 26.470 ;
        RECT 170.760 26.340 171.040 27.280 ;
        RECT 162.100 25.250 163.100 26.130 ;
        RECT 168.920 25.880 171.040 26.340 ;
        RECT 168.920 25.560 170.760 25.880 ;
        RECT 169.600 24.760 170.600 25.560 ;
        RECT 153.290 23.475 159.800 23.725 ;
        RECT 172.005 23.900 172.225 29.540 ;
        RECT 173.260 28.150 173.560 29.570 ;
        RECT 176.200 29.530 176.460 31.100 ;
        RECT 178.020 29.530 178.290 40.855 ;
        RECT 178.720 29.530 178.990 47.475 ;
        RECT 176.200 29.260 180.660 29.530 ;
        RECT 176.200 29.050 176.460 29.260 ;
        RECT 173.830 28.790 176.460 29.050 ;
        RECT 177.435 28.170 180.570 28.390 ;
        RECT 173.190 28.080 175.020 28.150 ;
        RECT 173.190 27.850 175.030 28.080 ;
        RECT 173.260 26.530 173.560 27.850 ;
        RECT 174.550 27.310 174.780 27.690 ;
        RECT 173.830 27.050 174.780 27.310 ;
        RECT 174.550 26.690 174.780 27.050 ;
        RECT 174.990 26.960 175.220 27.690 ;
        RECT 174.990 26.770 175.890 26.960 ;
        RECT 174.990 26.690 175.220 26.770 ;
        RECT 173.260 26.520 174.340 26.530 ;
        RECT 174.740 26.520 175.030 26.530 ;
        RECT 173.260 26.280 175.090 26.520 ;
        RECT 175.700 25.970 175.890 26.770 ;
        RECT 173.930 25.675 175.890 25.970 ;
        RECT 173.930 25.340 175.830 25.675 ;
        RECT 174.430 24.160 175.430 25.340 ;
        RECT 177.435 23.900 177.655 28.170 ;
        RECT 180.350 27.330 180.570 28.170 ;
        RECT 172.005 23.680 177.655 23.900 ;
        RECT 88.350 22.200 155.380 22.520 ;
        RECT 14.890 18.750 15.150 19.070 ;
        RECT 18.260 19.025 18.490 19.230 ;
        RECT 18.730 19.025 18.960 19.230 ;
        RECT 19.300 18.220 19.530 19.230 ;
        RECT 14.860 17.080 15.180 17.340 ;
        RECT 14.920 16.750 15.120 17.080 ;
        RECT 47.300 17.070 47.740 21.820 ;
        RECT 2.210 16.705 15.280 16.750 ;
        RECT -1.945 16.395 15.280 16.705 ;
        RECT -1.945 3.470 -1.635 16.395 ;
        RECT 2.210 16.230 15.280 16.395 ;
        RECT 37.840 16.630 47.740 17.070 ;
        RECT 114.940 20.195 120.590 20.415 ;
        RECT 23.490 13.800 23.720 13.900 ;
        RECT 22.480 13.620 23.720 13.800 ;
        RECT 3.130 13.140 3.360 13.335 ;
        RECT 11.020 13.150 11.250 13.405 ;
        RECT 3.130 12.950 4.470 13.140 ;
        RECT 3.130 12.795 3.360 12.950 ;
        RECT 4.280 11.760 4.470 12.950 ;
        RECT 9.840 12.970 11.250 13.150 ;
        RECT 9.840 11.810 10.020 12.970 ;
        RECT 11.020 12.865 11.250 12.970 ;
        RECT 11.490 13.250 11.720 13.405 ;
        RECT 11.490 13.080 13.050 13.250 ;
        RECT 11.490 12.865 11.720 13.080 ;
        RECT 10.590 12.000 12.150 12.150 ;
        RECT 10.420 11.980 12.260 12.000 ;
        RECT 10.420 11.850 12.360 11.980 ;
        RECT 10.420 11.810 12.620 11.850 ;
        RECT 4.280 11.480 8.400 11.760 ;
        RECT 9.840 11.630 12.620 11.810 ;
        RECT 4.280 11.325 4.470 11.480 ;
        RECT 1.935 11.135 4.470 11.325 ;
        RECT 1.935 10.930 2.125 11.135 ;
        RECT 1.900 10.610 2.160 10.930 ;
        RECT 8.120 10.245 8.400 11.480 ;
        RECT 12.270 11.590 12.620 11.630 ;
        RECT 12.270 10.680 12.450 11.590 ;
        RECT 12.230 10.360 12.490 10.680 ;
        RECT 8.120 10.195 10.030 10.245 ;
        RECT 12.880 10.195 13.050 13.080 ;
        RECT 22.480 12.770 22.660 13.620 ;
        RECT 23.490 13.480 23.720 13.620 ;
        RECT 34.360 13.065 34.590 13.120 ;
        RECT 34.360 12.875 35.535 13.065 ;
        RECT 23.060 12.770 24.620 12.810 ;
        RECT 17.130 12.590 24.620 12.770 ;
        RECT 34.360 12.700 34.590 12.875 ;
        RECT 17.130 12.310 17.310 12.590 ;
        RECT 23.060 12.580 24.620 12.590 ;
        RECT 17.090 11.990 17.350 12.310 ;
        RECT 33.460 11.985 35.020 12.030 ;
        RECT 35.345 11.985 35.535 12.875 ;
        RECT 13.280 11.810 13.540 11.880 ;
        RECT 13.280 11.630 19.230 11.810 ;
        RECT 33.460 11.800 35.535 11.985 ;
        RECT 13.280 11.560 13.540 11.630 ;
        RECT 17.060 10.960 17.380 11.220 ;
        RECT 8.120 10.080 13.050 10.195 ;
        RECT 8.120 10.020 8.400 10.080 ;
        RECT 9.585 10.025 13.050 10.080 ;
        RECT 1.870 9.805 2.190 9.840 ;
        RECT 2.550 9.805 2.780 9.900 ;
        RECT 3.020 9.810 3.250 9.900 ;
        RECT 1.870 9.615 2.780 9.805 ;
        RECT 1.870 9.580 2.190 9.615 ;
        RECT 2.550 9.480 2.780 9.615 ;
        RECT 3.010 9.600 4.250 9.810 ;
        RECT 3.020 9.480 3.250 9.600 ;
        RECT 4.040 8.835 4.250 9.600 ;
        RECT 3.235 8.820 4.250 8.835 ;
        RECT 2.040 8.625 4.250 8.820 ;
        RECT 2.040 8.100 3.790 8.625 ;
        RECT 2.890 3.470 3.200 8.100 ;
        RECT 9.050 7.400 9.310 7.435 ;
        RECT 8.195 7.150 9.310 7.400 ;
        RECT 8.195 6.850 8.445 7.150 ;
        RECT 9.050 7.115 9.310 7.150 ;
        RECT 7.430 6.600 8.450 6.850 ;
        RECT 9.585 6.775 9.755 10.025 ;
        RECT 12.200 9.420 12.520 9.680 ;
        RECT 10.100 7.400 10.420 7.405 ;
        RECT 10.100 7.150 11.640 7.400 ;
        RECT 10.100 7.145 10.420 7.150 ;
        RECT 11.335 7.140 11.625 7.150 ;
        RECT 11.130 6.775 11.360 6.980 ;
        RECT 9.585 6.605 11.360 6.775 ;
        RECT 7.430 3.470 7.680 6.600 ;
        RECT 8.195 6.345 8.445 6.600 ;
        RECT 11.130 6.560 11.360 6.605 ;
        RECT 11.600 6.810 11.830 6.980 ;
        RECT 12.270 6.810 12.450 9.420 ;
        RECT 11.600 6.630 12.450 6.810 ;
        RECT 11.600 6.560 11.830 6.630 ;
        RECT 12.270 6.440 12.450 6.630 ;
        RECT 11.335 6.345 11.625 6.400 ;
        RECT 8.195 6.095 11.655 6.345 ;
        RECT 11.930 6.260 12.450 6.440 ;
        RECT 11.930 5.890 12.110 6.260 ;
        RECT 10.700 5.660 12.260 5.890 ;
        RECT 17.130 5.380 17.310 10.960 ;
        RECT 19.050 8.110 19.230 11.630 ;
        RECT 34.715 11.795 35.535 11.800 ;
        RECT 22.070 8.510 23.100 8.690 ;
        RECT 22.070 8.110 22.250 8.510 ;
        RECT 22.795 8.450 23.085 8.510 ;
        RECT 22.590 8.190 22.820 8.290 ;
        RECT 23.060 8.190 23.290 8.290 ;
        RECT 23.630 8.190 23.860 9.050 ;
        RECT 19.050 7.930 22.250 8.110 ;
        RECT 22.560 8.000 26.230 8.190 ;
        RECT 21.930 7.680 22.110 7.930 ;
        RECT 22.590 7.870 22.820 8.000 ;
        RECT 23.060 7.870 23.290 8.000 ;
        RECT 22.795 7.680 23.085 7.710 ;
        RECT 21.930 7.500 23.085 7.680 ;
        RECT 22.795 7.480 23.085 7.500 ;
        RECT 23.630 7.110 23.860 8.000 ;
        RECT 26.040 5.615 26.230 8.000 ;
        RECT 34.715 5.615 34.905 11.795 ;
        RECT 26.040 5.425 34.905 5.615 ;
        RECT 17.060 5.120 17.380 5.380 ;
        RECT 17.060 3.840 17.380 4.100 ;
        RECT -1.945 3.420 16.930 3.470 ;
        RECT 17.130 3.420 17.310 3.840 ;
        RECT -1.945 3.170 17.440 3.420 ;
        RECT -1.945 3.160 8.970 3.170 ;
        RECT 11.090 3.160 17.440 3.170 ;
        RECT 6.830 -4.750 7.270 3.160 ;
        RECT 13.605 0.840 13.915 3.160 ;
        RECT 26.040 2.450 26.230 5.425 ;
        RECT 26.005 2.130 26.265 2.450 ;
        RECT 25.975 0.960 26.295 1.220 ;
        RECT 13.605 0.495 14.280 0.840 ;
        RECT 13.700 -0.800 14.280 0.495 ;
        RECT 26.040 0.410 26.230 0.960 ;
        RECT 23.795 0.180 29.865 0.410 ;
        RECT 15.280 -0.060 15.480 -0.030 ;
        RECT 15.035 -0.290 21.105 -0.060 ;
        RECT 14.010 -1.160 14.210 -0.800 ;
        RECT 15.280 -1.160 15.480 -0.290 ;
        RECT 14.010 -1.360 15.480 -1.160 ;
        RECT 6.830 -4.780 37.490 -4.750 ;
        RECT 37.840 -4.780 38.280 16.630 ;
        RECT 112.220 15.925 113.220 16.440 ;
        RECT 114.940 15.925 115.160 20.195 ;
        RECT 117.165 18.755 118.165 19.935 ;
        RECT 116.765 18.420 118.665 18.755 ;
        RECT 116.705 18.125 118.665 18.420 ;
        RECT 116.705 17.325 116.895 18.125 ;
        RECT 117.505 17.575 119.335 17.815 ;
        RECT 117.565 17.565 117.855 17.575 ;
        RECT 118.255 17.565 119.335 17.575 ;
        RECT 117.375 17.325 117.605 17.405 ;
        RECT 116.705 17.135 117.605 17.325 ;
        RECT 117.375 16.405 117.605 17.135 ;
        RECT 117.815 17.045 118.045 17.405 ;
        RECT 117.815 16.785 118.765 17.045 ;
        RECT 117.815 16.405 118.045 16.785 ;
        RECT 119.035 16.245 119.335 17.565 ;
        RECT 117.565 16.015 119.405 16.245 ;
        RECT 117.575 15.945 119.405 16.015 ;
        RECT 112.220 15.705 115.160 15.925 ;
        RECT 112.220 15.440 113.220 15.705 ;
        RECT 116.135 15.045 118.765 15.305 ;
        RECT 116.135 14.835 116.395 15.045 ;
        RECT 111.935 14.565 116.395 14.835 ;
        RECT 52.060 13.405 52.330 13.415 ;
        RECT 59.660 13.405 59.930 13.455 ;
        RECT 67.310 13.405 67.580 13.415 ;
        RECT 75.150 13.405 75.420 13.455 ;
        RECT 83.070 13.405 83.340 13.415 ;
        RECT 90.740 13.405 91.010 13.425 ;
        RECT 50.850 13.135 98.310 13.405 ;
        RECT 48.350 11.890 48.580 11.935 ;
        RECT 50.290 11.890 50.610 11.905 ;
        RECT 48.350 11.660 50.610 11.890 ;
        RECT 48.350 11.255 48.580 11.660 ;
        RECT 50.290 11.645 50.610 11.660 ;
        RECT 47.920 9.665 48.920 11.255 ;
        RECT 48.170 9.035 48.410 9.665 ;
        RECT 46.000 9.025 48.410 9.035 ;
        RECT 45.530 8.835 48.410 9.025 ;
        RECT 45.530 8.795 47.090 8.835 ;
        RECT 44.580 8.515 46.480 8.525 ;
        RECT 44.570 8.265 46.480 8.515 ;
        RECT 44.570 6.095 44.800 8.265 ;
        RECT 45.960 7.895 46.190 7.995 ;
        RECT 48.170 7.895 48.410 8.835 ;
        RECT 45.960 7.655 48.410 7.895 ;
        RECT 45.960 7.205 46.190 7.655 ;
        RECT 46.430 6.575 46.660 7.155 ;
        RECT 46.430 6.445 47.620 6.575 ;
        RECT 50.850 6.450 51.120 13.135 ;
        RECT 52.060 9.995 52.330 13.135 ;
        RECT 52.720 11.890 52.980 11.935 ;
        RECT 54.550 11.890 55.550 12.175 ;
        RECT 58.850 11.890 59.170 11.905 ;
        RECT 52.720 11.660 59.170 11.890 ;
        RECT 52.720 11.615 52.980 11.660 ;
        RECT 54.550 11.445 55.550 11.660 ;
        RECT 58.850 11.645 59.170 11.660 ;
        RECT 53.670 11.125 53.990 11.135 ;
        RECT 54.240 11.125 55.970 11.445 ;
        RECT 53.670 10.885 55.970 11.125 ;
        RECT 53.670 10.875 53.990 10.885 ;
        RECT 54.240 10.565 55.970 10.885 ;
        RECT 54.925 10.215 55.215 10.265 ;
        RECT 53.440 10.065 55.215 10.215 ;
        RECT 51.780 9.635 52.780 9.995 ;
        RECT 53.450 9.635 53.640 10.065 ;
        RECT 54.925 10.035 55.215 10.065 ;
        RECT 59.660 10.045 59.930 13.135 ;
        RECT 60.410 11.890 60.670 11.935 ;
        RECT 62.140 11.890 63.140 12.225 ;
        RECT 66.670 11.890 66.990 11.905 ;
        RECT 60.410 11.660 66.990 11.890 ;
        RECT 60.410 11.615 60.670 11.660 ;
        RECT 62.140 11.495 63.140 11.660 ;
        RECT 66.670 11.645 66.990 11.660 ;
        RECT 61.260 11.175 61.580 11.185 ;
        RECT 61.830 11.175 63.560 11.495 ;
        RECT 61.260 10.935 63.560 11.175 ;
        RECT 61.260 10.925 61.580 10.935 ;
        RECT 61.830 10.615 63.560 10.935 ;
        RECT 62.515 10.265 62.805 10.315 ;
        RECT 61.030 10.115 62.805 10.265 ;
        RECT 51.780 9.365 53.640 9.635 ;
        RECT 51.780 8.995 52.780 9.365 ;
        RECT 53.450 8.865 53.640 9.365 ;
        RECT 53.970 9.615 54.230 9.655 ;
        RECT 54.720 9.615 54.950 9.830 ;
        RECT 53.970 9.375 54.950 9.615 ;
        RECT 53.970 9.335 54.230 9.375 ;
        RECT 54.720 9.110 54.950 9.375 ;
        RECT 55.190 9.775 55.420 9.830 ;
        RECT 55.620 9.775 55.940 9.820 ;
        RECT 55.190 9.605 55.940 9.775 ;
        RECT 55.190 9.110 55.420 9.605 ;
        RECT 55.620 9.560 55.940 9.605 ;
        RECT 59.370 9.685 60.370 10.045 ;
        RECT 61.040 9.685 61.230 10.115 ;
        RECT 62.515 10.085 62.805 10.115 ;
        RECT 67.310 10.065 67.580 13.135 ;
        RECT 67.850 11.890 68.110 11.935 ;
        RECT 69.750 11.890 70.750 12.245 ;
        RECT 74.650 11.890 74.910 11.935 ;
        RECT 67.850 11.660 74.910 11.890 ;
        RECT 67.850 11.615 68.110 11.660 ;
        RECT 69.750 11.515 70.750 11.660 ;
        RECT 74.650 11.615 74.910 11.660 ;
        RECT 68.870 11.195 69.190 11.205 ;
        RECT 69.440 11.195 71.170 11.515 ;
        RECT 68.870 10.955 71.170 11.195 ;
        RECT 68.870 10.945 69.190 10.955 ;
        RECT 69.440 10.635 71.170 10.955 ;
        RECT 70.125 10.285 70.415 10.335 ;
        RECT 68.640 10.135 70.415 10.285 ;
        RECT 59.370 9.415 61.230 9.685 ;
        RECT 59.370 9.045 60.370 9.415 ;
        RECT 61.040 8.915 61.230 9.415 ;
        RECT 61.560 9.665 61.820 9.705 ;
        RECT 62.310 9.665 62.540 9.880 ;
        RECT 61.560 9.425 62.540 9.665 ;
        RECT 61.560 9.385 61.820 9.425 ;
        RECT 62.310 9.160 62.540 9.425 ;
        RECT 62.780 9.825 63.010 9.880 ;
        RECT 63.210 9.825 63.530 9.870 ;
        RECT 62.780 9.655 63.530 9.825 ;
        RECT 62.780 9.160 63.010 9.655 ;
        RECT 63.210 9.610 63.530 9.655 ;
        RECT 66.980 9.705 67.980 10.065 ;
        RECT 68.650 9.705 68.840 10.135 ;
        RECT 70.125 10.105 70.415 10.135 ;
        RECT 75.150 10.025 75.420 13.135 ;
        RECT 75.770 11.890 76.030 11.935 ;
        RECT 77.750 11.890 78.750 12.205 ;
        RECT 82.260 11.890 82.580 11.905 ;
        RECT 75.770 11.660 82.580 11.890 ;
        RECT 75.770 11.615 76.030 11.660 ;
        RECT 77.750 11.475 78.750 11.660 ;
        RECT 82.260 11.645 82.580 11.660 ;
        RECT 76.870 11.155 77.190 11.165 ;
        RECT 77.440 11.155 79.170 11.475 ;
        RECT 76.870 10.915 79.170 11.155 ;
        RECT 76.870 10.905 77.190 10.915 ;
        RECT 77.440 10.595 79.170 10.915 ;
        RECT 78.125 10.245 78.415 10.295 ;
        RECT 76.640 10.095 78.415 10.245 ;
        RECT 66.980 9.435 68.840 9.705 ;
        RECT 66.980 9.065 67.980 9.435 ;
        RECT 67.310 9.005 67.580 9.065 ;
        RECT 62.515 8.915 62.805 8.955 ;
        RECT 68.650 8.935 68.840 9.435 ;
        RECT 69.170 9.685 69.430 9.725 ;
        RECT 69.920 9.685 70.150 9.900 ;
        RECT 69.170 9.445 70.150 9.685 ;
        RECT 69.170 9.405 69.430 9.445 ;
        RECT 69.920 9.180 70.150 9.445 ;
        RECT 70.390 9.845 70.620 9.900 ;
        RECT 70.820 9.845 71.140 9.890 ;
        RECT 70.390 9.675 71.140 9.845 ;
        RECT 70.390 9.180 70.620 9.675 ;
        RECT 70.820 9.630 71.140 9.675 ;
        RECT 74.980 9.665 75.980 10.025 ;
        RECT 76.650 9.665 76.840 10.095 ;
        RECT 78.125 10.065 78.415 10.095 ;
        RECT 83.070 10.045 83.340 13.135 ;
        RECT 83.640 11.890 83.900 11.935 ;
        RECT 85.560 11.890 86.560 12.225 ;
        RECT 90.190 11.890 90.510 11.905 ;
        RECT 83.640 11.660 90.510 11.890 ;
        RECT 83.640 11.615 83.900 11.660 ;
        RECT 85.560 11.495 86.560 11.660 ;
        RECT 90.190 11.645 90.510 11.660 ;
        RECT 84.680 11.175 85.000 11.185 ;
        RECT 85.250 11.175 86.980 11.495 ;
        RECT 84.680 10.935 86.980 11.175 ;
        RECT 84.680 10.925 85.000 10.935 ;
        RECT 85.250 10.615 86.980 10.935 ;
        RECT 85.935 10.265 86.225 10.315 ;
        RECT 84.450 10.115 86.225 10.265 ;
        RECT 74.980 9.395 76.840 9.665 ;
        RECT 74.980 9.025 75.980 9.395 ;
        RECT 70.125 8.935 70.415 8.975 ;
        RECT 54.925 8.865 55.215 8.905 ;
        RECT 53.450 8.715 55.240 8.865 ;
        RECT 61.040 8.765 62.830 8.915 ;
        RECT 68.650 8.785 70.440 8.935 ;
        RECT 76.650 8.895 76.840 9.395 ;
        RECT 77.170 9.645 77.430 9.685 ;
        RECT 77.920 9.645 78.150 9.860 ;
        RECT 77.170 9.405 78.150 9.645 ;
        RECT 77.170 9.365 77.430 9.405 ;
        RECT 77.920 9.140 78.150 9.405 ;
        RECT 78.390 9.805 78.620 9.860 ;
        RECT 78.820 9.805 79.140 9.850 ;
        RECT 78.390 9.635 79.140 9.805 ;
        RECT 78.390 9.140 78.620 9.635 ;
        RECT 78.820 9.590 79.140 9.635 ;
        RECT 82.790 9.685 83.790 10.045 ;
        RECT 84.460 9.685 84.650 10.115 ;
        RECT 85.935 10.085 86.225 10.115 ;
        RECT 90.740 10.025 91.010 13.135 ;
        RECT 91.400 11.890 91.660 11.935 ;
        RECT 93.150 11.890 94.150 12.205 ;
        RECT 97.420 11.890 97.740 11.905 ;
        RECT 91.400 11.660 97.740 11.890 ;
        RECT 91.400 11.615 91.660 11.660 ;
        RECT 93.150 11.475 94.150 11.660 ;
        RECT 97.420 11.645 97.740 11.660 ;
        RECT 92.270 11.155 92.590 11.165 ;
        RECT 92.840 11.155 94.570 11.475 ;
        RECT 92.270 10.915 94.570 11.155 ;
        RECT 92.270 10.905 92.590 10.915 ;
        RECT 92.840 10.595 94.570 10.915 ;
        RECT 93.525 10.245 93.815 10.295 ;
        RECT 92.040 10.095 93.815 10.245 ;
        RECT 82.790 9.415 84.650 9.685 ;
        RECT 82.790 9.045 83.790 9.415 ;
        RECT 83.070 9.005 83.340 9.045 ;
        RECT 78.125 8.895 78.415 8.935 ;
        RECT 84.460 8.915 84.650 9.415 ;
        RECT 84.980 9.665 85.240 9.705 ;
        RECT 85.730 9.665 85.960 9.880 ;
        RECT 84.980 9.425 85.960 9.665 ;
        RECT 84.980 9.385 85.240 9.425 ;
        RECT 85.730 9.160 85.960 9.425 ;
        RECT 86.200 9.825 86.430 9.880 ;
        RECT 86.630 9.825 86.950 9.870 ;
        RECT 86.200 9.655 86.950 9.825 ;
        RECT 86.200 9.160 86.430 9.655 ;
        RECT 86.630 9.610 86.950 9.655 ;
        RECT 90.380 9.665 91.380 10.025 ;
        RECT 92.050 9.665 92.240 10.095 ;
        RECT 93.525 10.065 93.815 10.095 ;
        RECT 98.040 9.995 98.310 13.135 ;
        RECT 98.500 11.890 98.760 11.935 ;
        RECT 100.540 11.890 101.540 12.175 ;
        RECT 98.500 11.885 101.540 11.890 ;
        RECT 98.500 11.660 107.605 11.885 ;
        RECT 98.500 11.615 98.760 11.660 ;
        RECT 100.540 11.635 107.605 11.660 ;
        RECT 100.540 11.445 101.540 11.635 ;
        RECT 99.660 11.125 99.980 11.135 ;
        RECT 100.230 11.125 101.960 11.445 ;
        RECT 99.660 10.885 101.960 11.125 ;
        RECT 99.660 10.875 99.980 10.885 ;
        RECT 100.230 10.565 101.960 10.885 ;
        RECT 100.915 10.215 101.205 10.265 ;
        RECT 99.430 10.065 101.205 10.215 ;
        RECT 90.380 9.395 92.240 9.665 ;
        RECT 90.380 9.025 91.380 9.395 ;
        RECT 90.740 9.015 91.010 9.025 ;
        RECT 85.935 8.915 86.225 8.955 ;
        RECT 62.515 8.725 62.805 8.765 ;
        RECT 70.125 8.745 70.415 8.785 ;
        RECT 76.650 8.745 78.440 8.895 ;
        RECT 84.460 8.765 86.250 8.915 ;
        RECT 92.050 8.895 92.240 9.395 ;
        RECT 92.570 9.645 92.830 9.685 ;
        RECT 93.320 9.645 93.550 9.860 ;
        RECT 92.570 9.405 93.550 9.645 ;
        RECT 92.570 9.365 92.830 9.405 ;
        RECT 93.320 9.140 93.550 9.405 ;
        RECT 93.790 9.805 94.020 9.860 ;
        RECT 94.220 9.805 94.540 9.850 ;
        RECT 93.790 9.635 94.540 9.805 ;
        RECT 93.790 9.140 94.020 9.635 ;
        RECT 94.220 9.590 94.540 9.635 ;
        RECT 97.770 9.635 98.770 9.995 ;
        RECT 99.440 9.635 99.630 10.065 ;
        RECT 100.915 10.035 101.205 10.065 ;
        RECT 107.355 9.945 107.605 11.635 ;
        RECT 97.770 9.365 99.630 9.635 ;
        RECT 97.770 8.995 98.770 9.365 ;
        RECT 93.525 8.895 93.815 8.935 ;
        RECT 54.925 8.675 55.215 8.715 ;
        RECT 78.125 8.705 78.415 8.745 ;
        RECT 85.935 8.725 86.225 8.765 ;
        RECT 92.050 8.745 93.840 8.895 ;
        RECT 99.440 8.865 99.630 9.365 ;
        RECT 99.960 9.615 100.220 9.655 ;
        RECT 100.710 9.615 100.940 9.830 ;
        RECT 99.960 9.375 100.940 9.615 ;
        RECT 99.960 9.335 100.220 9.375 ;
        RECT 100.710 9.110 100.940 9.375 ;
        RECT 101.180 9.775 101.410 9.830 ;
        RECT 101.610 9.775 101.930 9.820 ;
        RECT 101.180 9.605 101.930 9.775 ;
        RECT 101.180 9.110 101.410 9.605 ;
        RECT 101.610 9.560 101.930 9.605 ;
        RECT 107.080 9.215 108.080 9.945 ;
        RECT 106.200 8.935 106.520 8.975 ;
        RECT 106.720 8.935 108.450 9.215 ;
        RECT 100.915 8.865 101.205 8.905 ;
        RECT 93.525 8.705 93.815 8.745 ;
        RECT 99.440 8.715 101.230 8.865 ;
        RECT 106.200 8.755 108.450 8.935 ;
        RECT 106.200 8.715 106.520 8.755 ;
        RECT 100.915 8.675 101.205 8.715 ;
        RECT 106.720 8.445 108.450 8.755 ;
        RECT 107.435 8.105 107.725 8.135 ;
        RECT 105.600 7.915 107.740 8.105 ;
        RECT 70.125 7.505 70.415 7.515 ;
        RECT 105.610 7.505 105.790 7.915 ;
        RECT 107.435 7.905 107.725 7.915 ;
        RECT 62.515 7.485 62.805 7.495 ;
        RECT 54.925 7.435 55.215 7.445 ;
        RECT 52.740 7.195 55.220 7.435 ;
        RECT 60.330 7.245 62.810 7.485 ;
        RECT 67.940 7.265 70.420 7.505 ;
        RECT 85.935 7.485 86.225 7.495 ;
        RECT 78.125 7.465 78.415 7.475 ;
        RECT 52.770 6.755 52.990 7.195 ;
        RECT 48.080 6.445 51.120 6.450 ;
        RECT 46.430 6.375 51.120 6.445 ;
        RECT 46.430 6.365 46.660 6.375 ;
        RECT 47.380 6.180 51.120 6.375 ;
        RECT 52.340 6.475 53.000 6.755 ;
        RECT 54.260 6.735 54.580 6.795 ;
        RECT 54.720 6.735 54.950 7.010 ;
        RECT 54.260 6.595 54.950 6.735 ;
        RECT 54.260 6.535 54.580 6.595 ;
        RECT 44.570 5.835 46.480 6.095 ;
        RECT 44.570 4.950 44.800 5.835 ;
        RECT 47.380 4.950 47.590 6.180 ;
        RECT 44.570 4.720 47.590 4.950 ;
        RECT 45.310 4.390 45.630 4.415 ;
        RECT 47.380 4.390 47.590 4.720 ;
        RECT 51.140 5.375 52.140 5.675 ;
        RECT 52.340 5.375 52.620 6.475 ;
        RECT 52.770 6.075 52.990 6.475 ;
        RECT 54.720 6.290 54.950 6.595 ;
        RECT 55.190 6.505 55.420 7.010 ;
        RECT 60.360 6.805 60.580 7.245 ;
        RECT 59.930 6.525 60.590 6.805 ;
        RECT 61.850 6.785 62.170 6.845 ;
        RECT 62.310 6.785 62.540 7.060 ;
        RECT 61.850 6.645 62.540 6.785 ;
        RECT 61.850 6.585 62.170 6.645 ;
        RECT 56.190 6.505 56.370 6.510 ;
        RECT 55.190 6.335 56.380 6.505 ;
        RECT 55.190 6.290 55.420 6.335 ;
        RECT 54.925 6.075 55.215 6.085 ;
        RECT 52.770 5.835 55.250 6.075 ;
        RECT 56.190 5.545 56.370 6.335 ;
        RECT 57.030 5.545 58.030 5.945 ;
        RECT 51.140 5.095 52.620 5.375 ;
        RECT 56.180 5.525 58.030 5.545 ;
        RECT 58.730 5.525 59.730 5.725 ;
        RECT 56.180 5.425 59.730 5.525 ;
        RECT 59.930 5.425 60.210 6.525 ;
        RECT 60.360 6.125 60.580 6.525 ;
        RECT 62.310 6.340 62.540 6.645 ;
        RECT 62.780 6.555 63.010 7.060 ;
        RECT 67.970 6.825 68.190 7.265 ;
        RECT 75.940 7.225 78.420 7.465 ;
        RECT 83.750 7.245 86.230 7.485 ;
        RECT 93.525 7.465 93.815 7.475 ;
        RECT 63.780 6.555 63.960 6.560 ;
        RECT 62.780 6.385 63.970 6.555 ;
        RECT 67.540 6.545 68.200 6.825 ;
        RECT 69.460 6.805 69.780 6.865 ;
        RECT 69.920 6.805 70.150 7.080 ;
        RECT 69.460 6.665 70.150 6.805 ;
        RECT 69.460 6.605 69.780 6.665 ;
        RECT 62.780 6.340 63.010 6.385 ;
        RECT 62.515 6.125 62.805 6.135 ;
        RECT 60.360 5.885 62.840 6.125 ;
        RECT 63.780 5.595 63.960 6.385 ;
        RECT 64.620 5.665 65.620 5.995 ;
        RECT 66.340 5.665 67.340 5.745 ;
        RECT 64.620 5.595 67.340 5.665 ;
        RECT 56.180 5.325 60.210 5.425 ;
        RECT 63.770 5.445 67.340 5.595 ;
        RECT 67.540 5.445 67.820 6.545 ;
        RECT 67.970 6.145 68.190 6.545 ;
        RECT 69.920 6.360 70.150 6.665 ;
        RECT 70.390 6.575 70.620 7.080 ;
        RECT 75.970 6.785 76.190 7.225 ;
        RECT 71.390 6.575 71.570 6.580 ;
        RECT 70.390 6.405 71.580 6.575 ;
        RECT 75.540 6.505 76.200 6.785 ;
        RECT 77.460 6.765 77.780 6.825 ;
        RECT 77.920 6.765 78.150 7.040 ;
        RECT 77.460 6.625 78.150 6.765 ;
        RECT 77.460 6.565 77.780 6.625 ;
        RECT 70.390 6.360 70.620 6.405 ;
        RECT 70.125 6.145 70.415 6.155 ;
        RECT 67.970 5.905 70.450 6.145 ;
        RECT 71.390 5.615 71.570 6.405 ;
        RECT 72.230 5.665 73.230 6.015 ;
        RECT 74.340 5.665 75.340 5.705 ;
        RECT 72.230 5.615 75.340 5.665 ;
        RECT 63.770 5.375 67.820 5.445 ;
        RECT 71.380 5.405 75.340 5.615 ;
        RECT 75.540 5.405 75.820 6.505 ;
        RECT 75.970 6.105 76.190 6.505 ;
        RECT 77.920 6.320 78.150 6.625 ;
        RECT 78.390 6.535 78.620 7.040 ;
        RECT 83.780 6.805 84.000 7.245 ;
        RECT 91.340 7.225 93.820 7.465 ;
        RECT 100.915 7.435 101.205 7.445 ;
        RECT 79.390 6.535 79.570 6.540 ;
        RECT 78.390 6.365 79.580 6.535 ;
        RECT 83.350 6.525 84.010 6.805 ;
        RECT 85.270 6.785 85.590 6.845 ;
        RECT 85.730 6.785 85.960 7.060 ;
        RECT 85.270 6.645 85.960 6.785 ;
        RECT 85.270 6.585 85.590 6.645 ;
        RECT 78.390 6.320 78.620 6.365 ;
        RECT 78.125 6.105 78.415 6.115 ;
        RECT 75.970 5.865 78.450 6.105 ;
        RECT 79.390 5.575 79.570 6.365 ;
        RECT 80.230 5.625 81.230 5.975 ;
        RECT 82.150 5.625 83.150 5.725 ;
        RECT 80.230 5.575 83.150 5.625 ;
        RECT 71.380 5.395 75.820 5.405 ;
        RECT 51.140 4.675 52.140 5.095 ;
        RECT 45.310 4.180 47.590 4.390 ;
        RECT 45.310 4.155 45.630 4.180 ;
        RECT 51.425 3.960 51.695 4.675 ;
        RECT 49.515 3.690 51.695 3.960 ;
        RECT 52.330 3.945 52.610 5.095 ;
        RECT 53.970 4.825 54.290 4.865 ;
        RECT 56.190 4.825 56.370 5.325 ;
        RECT 57.030 5.165 60.210 5.325 ;
        RECT 57.030 4.945 58.030 5.165 ;
        RECT 58.730 5.145 60.210 5.165 ;
        RECT 53.970 4.645 56.370 4.825 ;
        RECT 58.730 4.725 59.730 5.145 ;
        RECT 53.970 4.605 54.290 4.645 ;
        RECT 56.190 4.625 56.370 4.645 ;
        RECT 52.770 4.075 55.250 4.315 ;
        RECT 52.770 3.945 52.960 4.075 ;
        RECT 54.935 4.065 55.225 4.075 ;
        RECT 41.300 3.025 42.300 3.445 ;
        RECT 44.620 3.435 46.460 3.665 ;
        RECT 44.640 3.120 44.840 3.435 ;
        RECT 46.155 3.425 46.445 3.435 ;
        RECT 44.105 3.025 44.840 3.120 ;
        RECT 41.300 2.850 44.840 3.025 ;
        RECT 45.310 3.180 45.630 3.205 ;
        RECT 45.950 3.180 46.180 3.265 ;
        RECT 45.310 2.970 46.180 3.180 ;
        RECT 45.310 2.945 45.630 2.970 ;
        RECT 41.300 2.755 44.375 2.850 ;
        RECT 41.300 2.445 42.300 2.755 ;
        RECT 44.105 -1.595 44.375 2.755 ;
        RECT 44.640 2.695 44.840 2.850 ;
        RECT 45.950 2.845 46.180 2.970 ;
        RECT 46.420 3.115 46.650 3.265 ;
        RECT 46.420 2.895 47.670 3.115 ;
        RECT 46.420 2.845 46.650 2.895 ;
        RECT 44.630 2.465 46.470 2.695 ;
        RECT 46.155 2.455 46.445 2.465 ;
        RECT 45.520 2.095 47.080 2.175 ;
        RECT 45.490 1.805 47.100 2.095 ;
        RECT 47.450 1.805 47.670 2.895 ;
        RECT 45.490 1.585 47.670 1.805 ;
        RECT 45.490 1.225 47.100 1.585 ;
        RECT 45.770 0.595 46.770 1.225 ;
        RECT 46.350 -0.385 46.590 0.595 ;
        RECT 48.940 -0.385 49.260 -0.375 ;
        RECT 46.350 -0.625 49.260 -0.385 ;
        RECT 48.940 -0.635 49.260 -0.625 ;
        RECT 48.015 -1.595 48.285 -1.565 ;
        RECT 44.105 -1.865 48.285 -1.595 ;
        RECT 48.015 -1.895 48.285 -1.865 ;
        RECT 49.515 -2.350 49.785 3.690 ;
        RECT 52.330 3.665 52.960 3.945 ;
        RECT 59.920 3.995 60.200 5.145 ;
        RECT 61.560 4.875 61.880 4.915 ;
        RECT 63.780 4.875 63.960 5.375 ;
        RECT 64.620 5.305 67.820 5.375 ;
        RECT 64.620 4.995 65.620 5.305 ;
        RECT 66.340 5.165 67.820 5.305 ;
        RECT 61.560 4.695 63.960 4.875 ;
        RECT 66.340 4.745 67.340 5.165 ;
        RECT 61.560 4.655 61.880 4.695 ;
        RECT 63.780 4.675 63.960 4.695 ;
        RECT 60.360 4.125 62.840 4.365 ;
        RECT 60.360 3.995 60.550 4.125 ;
        RECT 62.525 4.115 62.815 4.125 ;
        RECT 52.770 3.335 52.960 3.665 ;
        RECT 54.000 3.835 54.260 3.905 ;
        RECT 54.730 3.835 54.960 3.905 ;
        RECT 54.000 3.655 54.960 3.835 ;
        RECT 54.000 3.585 54.260 3.655 ;
        RECT 54.580 3.645 54.960 3.655 ;
        RECT 54.730 3.485 54.960 3.645 ;
        RECT 55.200 3.715 55.430 3.905 ;
        RECT 59.920 3.715 60.550 3.995 ;
        RECT 67.530 4.015 67.810 5.165 ;
        RECT 69.170 4.895 69.490 4.935 ;
        RECT 71.390 4.895 71.570 5.395 ;
        RECT 72.230 5.305 75.820 5.395 ;
        RECT 79.380 5.425 83.150 5.575 ;
        RECT 83.350 5.425 83.630 6.525 ;
        RECT 83.780 6.125 84.000 6.525 ;
        RECT 85.730 6.340 85.960 6.645 ;
        RECT 86.200 6.555 86.430 7.060 ;
        RECT 91.370 6.785 91.590 7.225 ;
        RECT 98.730 7.195 101.210 7.435 ;
        RECT 105.010 7.255 105.790 7.505 ;
        RECT 87.200 6.555 87.380 6.560 ;
        RECT 86.200 6.385 87.390 6.555 ;
        RECT 90.940 6.505 91.600 6.785 ;
        RECT 92.860 6.765 93.180 6.825 ;
        RECT 93.320 6.765 93.550 7.040 ;
        RECT 92.860 6.625 93.550 6.765 ;
        RECT 92.860 6.565 93.180 6.625 ;
        RECT 86.200 6.340 86.430 6.385 ;
        RECT 85.935 6.125 86.225 6.135 ;
        RECT 83.780 5.885 86.260 6.125 ;
        RECT 87.200 5.595 87.380 6.385 ;
        RECT 88.040 5.625 89.040 5.995 ;
        RECT 89.740 5.625 90.740 5.705 ;
        RECT 88.040 5.595 90.740 5.625 ;
        RECT 79.380 5.355 83.630 5.425 ;
        RECT 87.190 5.405 90.740 5.595 ;
        RECT 90.940 5.405 91.220 6.505 ;
        RECT 91.370 6.105 91.590 6.505 ;
        RECT 93.320 6.320 93.550 6.625 ;
        RECT 93.790 6.535 94.020 7.040 ;
        RECT 98.760 6.755 98.980 7.195 ;
        RECT 94.790 6.535 94.970 6.540 ;
        RECT 93.790 6.365 94.980 6.535 ;
        RECT 98.330 6.475 98.990 6.755 ;
        RECT 100.250 6.735 100.570 6.795 ;
        RECT 100.710 6.735 100.940 7.010 ;
        RECT 100.250 6.595 100.940 6.735 ;
        RECT 100.250 6.535 100.570 6.595 ;
        RECT 93.790 6.320 94.020 6.365 ;
        RECT 93.525 6.105 93.815 6.115 ;
        RECT 91.370 5.865 93.850 6.105 ;
        RECT 94.790 5.575 94.970 6.365 ;
        RECT 95.630 5.575 96.630 5.975 ;
        RECT 97.130 5.575 98.130 5.675 ;
        RECT 87.190 5.375 91.220 5.405 ;
        RECT 72.230 5.015 73.230 5.305 ;
        RECT 74.340 5.125 75.820 5.305 ;
        RECT 69.170 4.715 71.570 4.895 ;
        RECT 69.170 4.675 69.490 4.715 ;
        RECT 71.390 4.695 71.570 4.715 ;
        RECT 74.340 4.705 75.340 5.125 ;
        RECT 67.970 4.145 70.450 4.385 ;
        RECT 67.970 4.015 68.160 4.145 ;
        RECT 70.135 4.135 70.425 4.145 ;
        RECT 55.200 3.545 56.380 3.715 ;
        RECT 55.200 3.485 55.430 3.545 ;
        RECT 52.770 3.095 55.250 3.335 ;
        RECT 54.070 2.190 54.390 2.235 ;
        RECT 56.205 2.190 56.375 3.545 ;
        RECT 60.360 3.385 60.550 3.715 ;
        RECT 61.590 3.885 61.850 3.955 ;
        RECT 62.320 3.885 62.550 3.955 ;
        RECT 61.590 3.705 62.550 3.885 ;
        RECT 61.590 3.635 61.850 3.705 ;
        RECT 62.170 3.695 62.550 3.705 ;
        RECT 62.320 3.535 62.550 3.695 ;
        RECT 62.790 3.765 63.020 3.955 ;
        RECT 62.790 3.595 63.970 3.765 ;
        RECT 67.530 3.735 68.160 4.015 ;
        RECT 75.530 3.975 75.810 5.125 ;
        RECT 77.170 4.855 77.490 4.895 ;
        RECT 79.390 4.855 79.570 5.355 ;
        RECT 80.230 5.265 83.630 5.355 ;
        RECT 80.230 4.975 81.230 5.265 ;
        RECT 82.150 5.145 83.630 5.265 ;
        RECT 77.170 4.675 79.570 4.855 ;
        RECT 82.150 4.725 83.150 5.145 ;
        RECT 77.170 4.635 77.490 4.675 ;
        RECT 79.390 4.655 79.570 4.675 ;
        RECT 75.970 4.105 78.450 4.345 ;
        RECT 75.970 3.975 76.160 4.105 ;
        RECT 78.135 4.095 78.425 4.105 ;
        RECT 62.790 3.535 63.020 3.595 ;
        RECT 60.360 3.145 62.840 3.385 ;
        RECT 54.070 2.020 56.375 2.190 ;
        RECT 61.660 2.240 61.980 2.285 ;
        RECT 63.795 2.240 63.965 3.595 ;
        RECT 67.970 3.405 68.160 3.735 ;
        RECT 69.200 3.905 69.460 3.975 ;
        RECT 69.930 3.905 70.160 3.975 ;
        RECT 69.200 3.725 70.160 3.905 ;
        RECT 69.200 3.655 69.460 3.725 ;
        RECT 69.780 3.715 70.160 3.725 ;
        RECT 69.930 3.555 70.160 3.715 ;
        RECT 70.400 3.785 70.630 3.975 ;
        RECT 70.400 3.615 71.580 3.785 ;
        RECT 75.530 3.695 76.160 3.975 ;
        RECT 83.340 3.995 83.620 5.145 ;
        RECT 84.980 4.875 85.300 4.915 ;
        RECT 87.200 4.875 87.380 5.375 ;
        RECT 88.040 5.265 91.220 5.375 ;
        RECT 94.780 5.375 98.130 5.575 ;
        RECT 98.330 5.375 98.610 6.475 ;
        RECT 98.760 6.075 98.980 6.475 ;
        RECT 100.710 6.290 100.940 6.595 ;
        RECT 101.180 6.505 101.410 7.010 ;
        RECT 102.180 6.505 102.360 6.510 ;
        RECT 101.180 6.335 102.370 6.505 ;
        RECT 101.180 6.290 101.410 6.335 ;
        RECT 100.915 6.075 101.205 6.085 ;
        RECT 98.760 5.835 101.240 6.075 ;
        RECT 102.180 5.545 102.360 6.335 ;
        RECT 103.020 5.625 104.020 5.945 ;
        RECT 105.020 5.625 105.190 7.255 ;
        RECT 105.610 6.765 105.790 7.255 ;
        RECT 106.230 7.455 106.490 7.525 ;
        RECT 107.230 7.455 107.460 7.700 ;
        RECT 106.230 7.275 107.460 7.455 ;
        RECT 106.230 7.205 106.490 7.275 ;
        RECT 107.230 6.980 107.460 7.275 ;
        RECT 107.700 7.445 107.930 7.700 ;
        RECT 107.700 7.255 108.900 7.445 ;
        RECT 107.700 6.980 107.930 7.255 ;
        RECT 107.435 6.765 107.725 6.775 ;
        RECT 105.610 6.575 107.750 6.765 ;
        RECT 107.435 6.545 107.725 6.575 ;
        RECT 103.020 5.545 105.190 5.625 ;
        RECT 94.780 5.355 98.610 5.375 ;
        RECT 88.040 4.995 89.040 5.265 ;
        RECT 89.740 5.125 91.220 5.265 ;
        RECT 84.980 4.695 87.380 4.875 ;
        RECT 89.740 4.705 90.740 5.125 ;
        RECT 84.980 4.655 85.300 4.695 ;
        RECT 87.200 4.675 87.380 4.695 ;
        RECT 83.780 4.125 86.260 4.365 ;
        RECT 83.780 3.995 83.970 4.125 ;
        RECT 85.945 4.115 86.235 4.125 ;
        RECT 70.400 3.555 70.630 3.615 ;
        RECT 67.970 3.165 70.450 3.405 ;
        RECT 61.660 2.070 63.965 2.240 ;
        RECT 69.270 2.260 69.590 2.305 ;
        RECT 71.405 2.260 71.575 3.615 ;
        RECT 75.970 3.365 76.160 3.695 ;
        RECT 77.200 3.865 77.460 3.935 ;
        RECT 77.930 3.865 78.160 3.935 ;
        RECT 77.200 3.685 78.160 3.865 ;
        RECT 77.200 3.615 77.460 3.685 ;
        RECT 77.780 3.675 78.160 3.685 ;
        RECT 77.930 3.515 78.160 3.675 ;
        RECT 78.400 3.745 78.630 3.935 ;
        RECT 78.400 3.575 79.580 3.745 ;
        RECT 83.340 3.715 83.970 3.995 ;
        RECT 90.930 3.975 91.210 5.125 ;
        RECT 92.570 4.855 92.890 4.895 ;
        RECT 94.790 4.855 94.970 5.355 ;
        RECT 95.630 5.215 98.610 5.355 ;
        RECT 102.170 5.355 105.190 5.545 ;
        RECT 108.705 6.155 108.895 7.255 ;
        RECT 109.360 6.155 110.360 6.645 ;
        RECT 108.705 5.895 110.360 6.155 ;
        RECT 102.170 5.325 104.020 5.355 ;
        RECT 95.630 4.975 96.630 5.215 ;
        RECT 97.130 5.095 98.610 5.215 ;
        RECT 92.570 4.675 94.970 4.855 ;
        RECT 97.130 4.675 98.130 5.095 ;
        RECT 92.570 4.635 92.890 4.675 ;
        RECT 94.790 4.655 94.970 4.675 ;
        RECT 91.370 4.105 93.850 4.345 ;
        RECT 91.370 3.975 91.560 4.105 ;
        RECT 93.535 4.095 93.825 4.105 ;
        RECT 78.400 3.515 78.630 3.575 ;
        RECT 75.970 3.125 78.450 3.365 ;
        RECT 69.270 2.090 71.575 2.260 ;
        RECT 77.270 2.220 77.590 2.265 ;
        RECT 79.405 2.220 79.575 3.575 ;
        RECT 83.780 3.385 83.970 3.715 ;
        RECT 85.010 3.885 85.270 3.955 ;
        RECT 85.740 3.885 85.970 3.955 ;
        RECT 85.010 3.705 85.970 3.885 ;
        RECT 85.010 3.635 85.270 3.705 ;
        RECT 85.590 3.695 85.970 3.705 ;
        RECT 85.740 3.535 85.970 3.695 ;
        RECT 86.210 3.765 86.440 3.955 ;
        RECT 86.210 3.595 87.390 3.765 ;
        RECT 90.930 3.695 91.560 3.975 ;
        RECT 98.320 3.945 98.600 5.095 ;
        RECT 99.960 4.825 100.280 4.865 ;
        RECT 102.180 4.825 102.360 5.325 ;
        RECT 103.020 4.945 104.020 5.325 ;
        RECT 99.960 4.645 102.360 4.825 ;
        RECT 99.960 4.605 100.280 4.645 ;
        RECT 102.180 4.625 102.360 4.645 ;
        RECT 98.760 4.075 101.240 4.315 ;
        RECT 98.760 3.945 98.950 4.075 ;
        RECT 100.925 4.065 101.215 4.075 ;
        RECT 86.210 3.535 86.440 3.595 ;
        RECT 83.780 3.145 86.260 3.385 ;
        RECT 61.660 2.025 61.980 2.070 ;
        RECT 69.270 2.045 69.590 2.090 ;
        RECT 77.270 2.050 79.575 2.220 ;
        RECT 85.080 2.240 85.400 2.285 ;
        RECT 87.215 2.240 87.385 3.595 ;
        RECT 91.370 3.365 91.560 3.695 ;
        RECT 92.600 3.865 92.860 3.935 ;
        RECT 93.330 3.865 93.560 3.935 ;
        RECT 92.600 3.685 93.560 3.865 ;
        RECT 92.600 3.615 92.860 3.685 ;
        RECT 93.180 3.675 93.560 3.685 ;
        RECT 93.330 3.515 93.560 3.675 ;
        RECT 93.800 3.745 94.030 3.935 ;
        RECT 93.800 3.575 94.980 3.745 ;
        RECT 98.320 3.665 98.950 3.945 ;
        RECT 93.800 3.515 94.030 3.575 ;
        RECT 91.370 3.125 93.850 3.365 ;
        RECT 85.080 2.070 87.385 2.240 ;
        RECT 92.670 2.220 92.990 2.265 ;
        RECT 94.805 2.220 94.975 3.575 ;
        RECT 98.760 3.335 98.950 3.665 ;
        RECT 99.990 3.835 100.250 3.905 ;
        RECT 100.720 3.835 100.950 3.905 ;
        RECT 99.990 3.655 100.950 3.835 ;
        RECT 99.990 3.585 100.250 3.655 ;
        RECT 100.570 3.645 100.950 3.655 ;
        RECT 100.720 3.485 100.950 3.645 ;
        RECT 101.190 3.715 101.420 3.905 ;
        RECT 101.190 3.545 102.370 3.715 ;
        RECT 101.190 3.485 101.420 3.545 ;
        RECT 98.760 3.095 101.240 3.335 ;
        RECT 54.070 1.975 54.390 2.020 ;
        RECT 77.270 2.005 77.590 2.050 ;
        RECT 85.080 2.025 85.400 2.070 ;
        RECT 92.670 2.050 94.975 2.220 ;
        RECT 100.060 2.190 100.380 2.235 ;
        RECT 102.195 2.190 102.365 3.545 ;
        RECT 92.670 2.005 92.990 2.050 ;
        RECT 100.060 2.020 102.365 2.190 ;
        RECT 100.060 1.975 100.380 2.020 ;
        RECT 62.535 1.885 62.825 1.915 ;
        RECT 70.145 1.905 70.435 1.935 ;
        RECT 54.945 1.835 55.235 1.865 ;
        RECT 52.090 1.545 53.090 1.775 ;
        RECT 53.390 1.615 55.250 1.835 ;
        RECT 53.390 1.545 53.610 1.615 ;
        RECT 52.090 1.325 53.610 1.545 ;
        RECT 59.680 1.595 60.680 1.825 ;
        RECT 60.980 1.665 62.840 1.885 ;
        RECT 60.980 1.595 61.200 1.665 ;
        RECT 54.070 1.350 54.390 1.395 ;
        RECT 54.740 1.350 54.970 1.475 ;
        RECT 52.090 0.775 53.090 1.325 ;
        RECT 53.380 0.895 53.600 1.325 ;
        RECT 54.070 1.180 54.970 1.350 ;
        RECT 54.070 1.135 54.390 1.180 ;
        RECT 54.650 1.150 54.970 1.180 ;
        RECT 54.740 1.055 54.970 1.150 ;
        RECT 55.210 1.295 55.440 1.475 ;
        RECT 59.680 1.375 61.200 1.595 ;
        RECT 67.290 1.615 68.290 1.845 ;
        RECT 68.590 1.685 70.450 1.905 ;
        RECT 78.145 1.865 78.435 1.895 ;
        RECT 85.955 1.885 86.245 1.915 ;
        RECT 68.590 1.615 68.810 1.685 ;
        RECT 61.660 1.400 61.980 1.445 ;
        RECT 62.330 1.400 62.560 1.525 ;
        RECT 55.210 1.125 55.940 1.295 ;
        RECT 55.210 1.055 55.440 1.125 ;
        RECT 50.190 -0.385 50.450 -0.345 ;
        RECT 51.800 -0.385 52.120 -0.375 ;
        RECT 50.190 -0.625 52.120 -0.385 ;
        RECT 50.190 -0.665 50.450 -0.625 ;
        RECT 51.800 -0.635 52.120 -0.625 ;
        RECT 52.340 -1.595 52.610 0.775 ;
        RECT 53.380 0.675 55.235 0.895 ;
        RECT 54.945 0.665 55.235 0.675 ;
        RECT 55.745 0.475 55.915 1.125 ;
        RECT 59.680 0.825 60.680 1.375 ;
        RECT 60.970 0.945 61.190 1.375 ;
        RECT 61.660 1.230 62.560 1.400 ;
        RECT 61.660 1.185 61.980 1.230 ;
        RECT 62.240 1.200 62.560 1.230 ;
        RECT 62.330 1.105 62.560 1.200 ;
        RECT 62.800 1.345 63.030 1.525 ;
        RECT 67.290 1.395 68.810 1.615 ;
        RECT 75.290 1.575 76.290 1.805 ;
        RECT 76.590 1.645 78.450 1.865 ;
        RECT 76.590 1.575 76.810 1.645 ;
        RECT 69.270 1.420 69.590 1.465 ;
        RECT 69.940 1.420 70.170 1.545 ;
        RECT 62.800 1.175 63.530 1.345 ;
        RECT 62.800 1.105 63.030 1.175 ;
        RECT 54.290 0.035 55.920 0.475 ;
        RECT 52.960 -0.385 53.220 -0.345 ;
        RECT 54.600 -0.385 55.600 0.035 ;
        RECT 59.370 -0.385 59.690 -0.375 ;
        RECT 52.960 -0.625 59.690 -0.385 ;
        RECT 52.960 -0.665 53.220 -0.625 ;
        RECT 54.600 -0.775 55.600 -0.625 ;
        RECT 59.370 -0.635 59.690 -0.625 ;
        RECT 59.940 -1.595 60.210 0.825 ;
        RECT 60.970 0.725 62.825 0.945 ;
        RECT 62.535 0.715 62.825 0.725 ;
        RECT 63.335 0.525 63.505 1.175 ;
        RECT 67.290 0.845 68.290 1.395 ;
        RECT 68.580 0.965 68.800 1.395 ;
        RECT 69.270 1.250 70.170 1.420 ;
        RECT 69.270 1.205 69.590 1.250 ;
        RECT 69.850 1.220 70.170 1.250 ;
        RECT 69.940 1.125 70.170 1.220 ;
        RECT 70.410 1.365 70.640 1.545 ;
        RECT 70.410 1.195 71.140 1.365 ;
        RECT 75.290 1.355 76.810 1.575 ;
        RECT 83.100 1.595 84.100 1.825 ;
        RECT 84.400 1.665 86.260 1.885 ;
        RECT 93.545 1.865 93.835 1.895 ;
        RECT 84.400 1.595 84.620 1.665 ;
        RECT 77.270 1.380 77.590 1.425 ;
        RECT 77.940 1.380 78.170 1.505 ;
        RECT 70.410 1.125 70.640 1.195 ;
        RECT 61.880 0.085 63.510 0.525 ;
        RECT 60.560 -0.385 60.820 -0.345 ;
        RECT 62.190 -0.385 63.190 0.085 ;
        RECT 66.980 -0.385 67.300 -0.375 ;
        RECT 60.560 -0.625 67.300 -0.385 ;
        RECT 60.560 -0.665 60.820 -0.625 ;
        RECT 62.190 -0.725 63.190 -0.625 ;
        RECT 66.980 -0.635 67.300 -0.625 ;
        RECT 67.620 -1.595 67.890 0.845 ;
        RECT 68.580 0.745 70.435 0.965 ;
        RECT 70.145 0.735 70.435 0.745 ;
        RECT 70.945 0.545 71.115 1.195 ;
        RECT 75.290 0.805 76.290 1.355 ;
        RECT 76.580 0.925 76.800 1.355 ;
        RECT 77.270 1.210 78.170 1.380 ;
        RECT 77.270 1.165 77.590 1.210 ;
        RECT 77.850 1.180 78.170 1.210 ;
        RECT 77.940 1.085 78.170 1.180 ;
        RECT 78.410 1.325 78.640 1.505 ;
        RECT 83.100 1.375 84.620 1.595 ;
        RECT 90.690 1.575 91.690 1.805 ;
        RECT 91.990 1.645 93.850 1.865 ;
        RECT 100.935 1.835 101.225 1.865 ;
        RECT 91.990 1.575 92.210 1.645 ;
        RECT 85.080 1.400 85.400 1.445 ;
        RECT 85.750 1.400 85.980 1.525 ;
        RECT 78.410 1.155 79.140 1.325 ;
        RECT 78.410 1.085 78.640 1.155 ;
        RECT 69.490 0.105 71.120 0.545 ;
        RECT 68.360 -0.385 68.620 -0.345 ;
        RECT 69.800 -0.385 70.800 0.105 ;
        RECT 74.860 -0.385 75.180 -0.375 ;
        RECT 68.360 -0.625 75.180 -0.385 ;
        RECT 68.360 -0.665 68.620 -0.625 ;
        RECT 69.800 -0.705 70.800 -0.625 ;
        RECT 74.860 -0.635 75.180 -0.625 ;
        RECT 75.500 -1.595 75.770 0.805 ;
        RECT 76.580 0.705 78.435 0.925 ;
        RECT 78.145 0.695 78.435 0.705 ;
        RECT 78.945 0.505 79.115 1.155 ;
        RECT 83.100 0.825 84.100 1.375 ;
        RECT 84.390 0.945 84.610 1.375 ;
        RECT 85.080 1.230 85.980 1.400 ;
        RECT 85.080 1.185 85.400 1.230 ;
        RECT 85.660 1.200 85.980 1.230 ;
        RECT 85.750 1.105 85.980 1.200 ;
        RECT 86.220 1.345 86.450 1.525 ;
        RECT 90.690 1.355 92.210 1.575 ;
        RECT 98.080 1.545 99.080 1.775 ;
        RECT 99.380 1.615 101.240 1.835 ;
        RECT 99.380 1.545 99.600 1.615 ;
        RECT 92.670 1.380 92.990 1.425 ;
        RECT 93.340 1.380 93.570 1.505 ;
        RECT 86.220 1.175 86.950 1.345 ;
        RECT 86.220 1.105 86.450 1.175 ;
        RECT 77.490 0.065 79.120 0.505 ;
        RECT 76.340 -0.385 76.600 -0.345 ;
        RECT 77.800 -0.385 78.800 0.065 ;
        RECT 82.730 -0.385 83.050 -0.375 ;
        RECT 76.340 -0.625 83.050 -0.385 ;
        RECT 76.340 -0.665 76.600 -0.625 ;
        RECT 77.800 -0.745 78.800 -0.625 ;
        RECT 82.730 -0.635 83.050 -0.625 ;
        RECT 83.450 -1.595 83.720 0.825 ;
        RECT 84.390 0.725 86.245 0.945 ;
        RECT 85.955 0.715 86.245 0.725 ;
        RECT 86.755 0.525 86.925 1.175 ;
        RECT 90.690 0.805 91.690 1.355 ;
        RECT 91.980 0.925 92.200 1.355 ;
        RECT 92.670 1.210 93.570 1.380 ;
        RECT 92.670 1.165 92.990 1.210 ;
        RECT 93.250 1.180 93.570 1.210 ;
        RECT 93.340 1.085 93.570 1.180 ;
        RECT 93.810 1.325 94.040 1.505 ;
        RECT 98.080 1.325 99.600 1.545 ;
        RECT 100.060 1.350 100.380 1.395 ;
        RECT 100.730 1.350 100.960 1.475 ;
        RECT 93.810 1.155 94.540 1.325 ;
        RECT 93.810 1.085 94.040 1.155 ;
        RECT 85.300 0.085 86.930 0.525 ;
        RECT 84.000 -0.385 84.260 -0.345 ;
        RECT 85.610 -0.385 86.610 0.085 ;
        RECT 90.670 -0.385 90.990 -0.375 ;
        RECT 84.000 -0.625 90.990 -0.385 ;
        RECT 84.000 -0.665 84.260 -0.625 ;
        RECT 85.610 -0.725 86.610 -0.625 ;
        RECT 90.670 -0.635 90.990 -0.625 ;
        RECT 91.170 -1.595 91.440 0.805 ;
        RECT 91.980 0.705 93.835 0.925 ;
        RECT 93.545 0.695 93.835 0.705 ;
        RECT 94.345 0.505 94.515 1.155 ;
        RECT 98.080 0.775 99.080 1.325 ;
        RECT 99.370 0.895 99.590 1.325 ;
        RECT 100.060 1.180 100.960 1.350 ;
        RECT 100.060 1.135 100.380 1.180 ;
        RECT 100.640 1.150 100.960 1.180 ;
        RECT 100.730 1.055 100.960 1.150 ;
        RECT 101.200 1.295 101.430 1.475 ;
        RECT 101.200 1.125 101.930 1.295 ;
        RECT 101.200 1.055 101.430 1.125 ;
        RECT 92.890 0.065 94.520 0.505 ;
        RECT 91.870 -0.385 92.130 -0.345 ;
        RECT 93.200 -0.385 94.200 0.065 ;
        RECT 97.920 -0.385 98.240 -0.375 ;
        RECT 91.870 -0.625 98.240 -0.385 ;
        RECT 91.870 -0.665 92.130 -0.625 ;
        RECT 93.200 -0.745 94.200 -0.625 ;
        RECT 97.920 -0.635 98.240 -0.625 ;
        RECT 98.590 -1.595 98.860 0.775 ;
        RECT 99.370 0.675 101.225 0.895 ;
        RECT 100.935 0.665 101.225 0.675 ;
        RECT 101.735 0.475 101.905 1.125 ;
        RECT 100.280 0.035 101.910 0.475 ;
        RECT 99.140 -0.385 99.400 -0.345 ;
        RECT 100.590 -0.385 101.590 0.035 ;
        RECT 103.540 -0.385 103.860 -0.375 ;
        RECT 99.140 -0.625 103.860 -0.385 ;
        RECT 99.140 -0.665 99.400 -0.625 ;
        RECT 100.590 -0.775 101.590 -0.625 ;
        RECT 103.540 -0.635 103.860 -0.625 ;
        RECT 50.645 -1.865 98.860 -1.595 ;
        RECT 52.340 -1.895 52.610 -1.865 ;
        RECT 83.450 -1.875 83.720 -1.865 ;
        RECT 91.170 -1.875 91.440 -1.865 ;
        RECT 104.215 -2.350 104.485 5.355 ;
        RECT 105.020 4.355 105.190 5.355 ;
        RECT 106.400 5.390 106.720 5.425 ;
        RECT 108.705 5.390 108.895 5.895 ;
        RECT 109.360 5.645 110.360 5.895 ;
        RECT 106.400 5.200 108.895 5.390 ;
        RECT 106.400 5.165 106.720 5.200 ;
        RECT 107.385 4.725 107.675 4.745 ;
        RECT 105.570 4.715 107.710 4.725 ;
        RECT 105.540 4.535 107.710 4.715 ;
        RECT 105.540 4.355 105.750 4.535 ;
        RECT 107.385 4.515 107.675 4.535 ;
        RECT 105.020 4.175 105.750 4.355 ;
        RECT 105.030 4.155 105.750 4.175 ;
        RECT 105.540 3.745 105.750 4.155 ;
        RECT 106.430 4.190 106.690 4.255 ;
        RECT 107.180 4.190 107.410 4.355 ;
        RECT 106.430 4.000 107.410 4.190 ;
        RECT 106.430 3.935 106.690 4.000 ;
        RECT 107.180 3.935 107.410 4.000 ;
        RECT 107.650 4.185 107.880 4.355 ;
        RECT 107.650 4.015 108.730 4.185 ;
        RECT 107.650 3.935 107.880 4.015 ;
        RECT 107.385 3.745 107.675 3.775 ;
        RECT 105.540 3.555 107.690 3.745 ;
        RECT 107.385 3.545 107.675 3.555 ;
        RECT 106.600 2.880 108.380 3.235 ;
        RECT 108.545 2.880 108.715 4.015 ;
        RECT 106.600 2.710 108.715 2.880 ;
        RECT 106.600 2.415 108.380 2.710 ;
        RECT 107.050 1.665 108.050 2.415 ;
        RECT 105.660 -0.385 105.920 -0.345 ;
        RECT 107.510 -0.385 107.750 1.665 ;
        RECT 105.660 -0.625 107.760 -0.385 ;
        RECT 105.660 -0.665 105.920 -0.625 ;
        RECT 49.515 -2.620 104.485 -2.350 ;
        RECT 113.605 -3.380 113.875 14.565 ;
        RECT 114.305 3.240 114.575 14.565 ;
        RECT 116.135 12.995 116.395 14.565 ;
        RECT 119.035 14.525 119.335 15.945 ;
        RECT 120.370 14.555 120.590 20.195 ;
        RECT 132.795 20.370 139.305 20.620 ;
        RECT 121.995 18.535 122.995 19.335 ;
        RECT 121.835 18.215 123.675 18.535 ;
        RECT 121.555 17.755 123.675 18.215 ;
        RECT 129.495 17.965 130.495 18.845 ;
        RECT 121.555 16.815 121.835 17.755 ;
        RECT 129.255 17.625 130.805 17.965 ;
        RECT 122.600 17.495 124.690 17.565 ;
        RECT 122.585 17.285 124.690 17.495 ;
        RECT 122.585 17.265 122.875 17.285 ;
        RECT 122.395 16.815 122.625 17.105 ;
        RECT 121.555 16.535 122.665 16.815 ;
        RECT 122.835 16.750 123.065 17.105 ;
        RECT 123.615 16.750 123.875 16.785 ;
        RECT 122.395 16.105 122.625 16.535 ;
        RECT 122.835 16.500 123.875 16.750 ;
        RECT 122.835 16.105 123.065 16.500 ;
        RECT 123.615 16.465 123.875 16.500 ;
        RECT 122.585 15.905 122.875 15.945 ;
        RECT 124.410 15.905 124.690 17.285 ;
        RECT 129.105 17.385 130.935 17.625 ;
        RECT 129.105 17.165 129.345 17.385 ;
        RECT 130.695 17.235 130.935 17.385 ;
        RECT 129.065 16.905 129.385 17.165 ;
        RECT 130.675 16.975 130.935 17.235 ;
        RECT 122.560 15.625 124.690 15.905 ;
        RECT 123.585 15.060 123.905 15.065 ;
        RECT 121.350 14.810 123.905 15.060 ;
        RECT 121.350 14.555 121.600 14.810 ;
        RECT 123.585 14.805 123.905 14.810 ;
        RECT 119.825 14.525 121.600 14.555 ;
        RECT 119.025 14.445 121.600 14.525 ;
        RECT 117.515 14.325 121.600 14.445 ;
        RECT 117.515 14.255 120.075 14.325 ;
        RECT 117.515 14.145 119.335 14.255 ;
        RECT 117.405 12.995 117.635 13.970 ;
        RECT 116.135 12.735 117.635 12.995 ;
        RECT 117.405 11.470 117.635 12.735 ;
        RECT 117.845 12.115 118.075 13.970 ;
        RECT 119.025 12.635 119.325 14.145 ;
        RECT 121.350 12.695 121.600 14.325 ;
        RECT 124.410 14.275 124.690 15.625 ;
        RECT 128.065 16.525 130.125 16.705 ;
        RECT 128.065 14.405 128.245 16.525 ;
        RECT 129.105 16.255 129.345 16.285 ;
        RECT 129.095 15.935 129.355 16.255 ;
        RECT 129.945 16.125 130.125 16.525 ;
        RECT 129.105 15.645 129.355 15.935 ;
        RECT 129.515 15.895 130.515 16.125 ;
        RECT 129.105 15.635 129.345 15.645 ;
        RECT 129.515 15.455 130.515 15.685 ;
        RECT 130.675 15.615 130.925 16.975 ;
        RECT 131.185 16.335 131.775 16.685 ;
        RECT 130.225 14.710 130.405 15.455 ;
        RECT 131.185 15.335 132.515 16.335 ;
        RECT 131.185 14.885 131.775 15.335 ;
        RECT 132.795 14.710 133.045 20.370 ;
        RECT 135.410 19.045 136.410 19.865 ;
        RECT 135.130 18.775 137.020 19.045 ;
        RECT 135.045 18.445 137.020 18.775 ;
        RECT 135.045 17.355 135.285 18.445 ;
        RECT 135.840 17.905 138.150 18.205 ;
        RECT 135.725 17.355 135.955 17.745 ;
        RECT 135.045 17.115 135.955 17.355 ;
        RECT 135.725 16.745 135.955 17.115 ;
        RECT 136.165 17.280 136.395 17.745 ;
        RECT 136.650 17.280 136.970 17.305 ;
        RECT 136.165 17.070 136.970 17.280 ;
        RECT 136.165 16.745 136.395 17.070 ;
        RECT 136.650 17.045 136.970 17.070 ;
        RECT 137.850 16.595 138.150 17.905 ;
        RECT 135.830 16.295 138.150 16.595 ;
        RECT 136.650 15.600 136.970 15.625 ;
        RECT 134.575 15.390 136.970 15.600 ;
        RECT 134.575 15.265 134.785 15.390 ;
        RECT 136.650 15.365 136.970 15.390 ;
        RECT 130.195 14.460 133.045 14.710 ;
        RECT 133.890 15.005 134.785 15.265 ;
        RECT 126.285 14.275 128.245 14.405 ;
        RECT 124.340 14.245 128.245 14.275 ;
        RECT 122.540 14.225 128.245 14.245 ;
        RECT 122.540 14.045 126.475 14.225 ;
        RECT 122.540 13.965 124.690 14.045 ;
        RECT 122.615 13.945 122.905 13.965 ;
        RECT 122.425 12.695 122.655 13.740 ;
        RECT 119.025 12.335 120.055 12.635 ;
        RECT 121.345 12.445 122.655 12.695 ;
        RECT 117.845 11.855 119.435 12.115 ;
        RECT 117.845 11.470 118.075 11.855 ;
        RECT 117.595 11.195 117.885 11.265 ;
        RECT 119.755 11.195 120.055 12.335 ;
        RECT 122.425 11.240 122.655 12.445 ;
        RECT 122.865 12.180 123.095 13.740 ;
        RECT 124.410 12.385 124.690 13.965 ;
        RECT 124.020 12.180 124.280 12.245 ;
        RECT 122.865 11.990 124.280 12.180 ;
        RECT 122.865 11.240 123.095 11.990 ;
        RECT 124.020 11.925 124.280 11.990 ;
        RECT 124.450 11.755 124.690 12.385 ;
        RECT 117.535 10.895 120.055 11.195 ;
        RECT 124.410 11.085 124.690 11.755 ;
        RECT 122.610 10.805 124.690 11.085 ;
        RECT 116.795 10.165 118.635 10.755 ;
        RECT 116.795 9.905 119.435 10.165 ;
        RECT 121.885 10.065 123.705 10.535 ;
        RECT 123.990 10.065 124.310 10.100 ;
        RECT 116.795 9.895 118.635 9.905 ;
        RECT 117.275 8.505 118.275 9.895 ;
        RECT 121.885 9.875 124.310 10.065 ;
        RECT 121.885 9.845 123.705 9.875 ;
        RECT 122.345 8.285 123.345 9.845 ;
        RECT 123.990 9.840 124.310 9.875 ;
        RECT 120.105 7.635 120.455 8.275 ;
        RECT 119.265 7.355 121.135 7.635 ;
        RECT 118.245 6.805 120.275 7.025 ;
        RECT 118.245 4.895 118.465 6.805 ;
        RECT 119.295 6.025 119.575 6.635 ;
        RECT 120.055 6.525 120.275 6.805 ;
        RECT 119.725 6.295 120.725 6.525 ;
        RECT 120.890 6.335 121.095 7.355 ;
        RECT 121.335 6.645 121.745 7.065 ;
        RECT 119.725 5.855 120.725 6.085 ;
        RECT 120.885 6.045 121.115 6.335 ;
        RECT 120.890 5.995 121.095 6.045 ;
        RECT 115.855 4.675 118.465 4.895 ;
        RECT 120.115 4.825 120.315 5.855 ;
        RECT 121.335 5.645 122.675 6.645 ;
        RECT 121.335 5.305 121.745 5.645 ;
        RECT 125.270 4.825 125.470 14.045 ;
        RECT 126.285 11.855 126.465 14.045 ;
        RECT 127.205 13.445 128.065 13.875 ;
        RECT 126.625 12.445 128.065 13.445 ;
        RECT 130.225 13.365 130.405 14.460 ;
        RECT 128.335 12.615 128.635 13.175 ;
        RECT 128.810 13.135 131.310 13.365 ;
        RECT 128.810 12.695 131.310 12.925 ;
        RECT 127.205 12.165 128.065 12.445 ;
        RECT 128.875 11.855 129.055 12.695 ;
        RECT 126.285 11.675 129.055 11.855 ;
        RECT 131.455 11.345 131.755 13.205 ;
        RECT 128.305 11.045 131.755 11.345 ;
        RECT 130.045 10.405 130.355 11.045 ;
        RECT 115.855 3.240 116.075 4.675 ;
        RECT 120.115 4.625 125.470 4.825 ;
        RECT 117.255 3.775 118.055 4.055 ;
        RECT 114.305 2.970 116.075 3.240 ;
        RECT 115.855 2.145 116.075 2.970 ;
        RECT 116.395 2.775 118.055 3.775 ;
        RECT 120.115 3.655 120.315 4.625 ;
        RECT 118.415 2.815 118.705 3.495 ;
        RECT 118.850 3.425 121.350 3.655 ;
        RECT 121.590 3.465 121.880 3.510 ;
        RECT 118.850 2.985 121.350 3.215 ;
        RECT 121.555 3.175 121.880 3.465 ;
        RECT 117.255 2.355 118.055 2.775 ;
        RECT 119.235 2.145 119.455 2.985 ;
        RECT 115.855 1.925 119.455 2.145 ;
        RECT 121.590 1.390 121.880 3.175 ;
        RECT 133.890 2.745 134.150 15.005 ;
        RECT 134.575 13.315 134.785 15.005 ;
        RECT 137.850 15.045 138.150 16.295 ;
        RECT 139.055 15.275 139.305 20.370 ;
        RECT 155.060 19.815 155.380 22.200 ;
        RECT 141.045 18.705 142.045 19.445 ;
        RECT 154.620 18.825 155.620 19.815 ;
        RECT 140.615 18.245 142.375 18.705 ;
        RECT 154.220 18.565 156.000 18.825 ;
        RECT 140.605 18.045 142.375 18.245 ;
        RECT 140.605 16.955 140.805 18.045 ;
        RECT 148.910 17.860 149.170 17.925 ;
        RECT 149.695 17.860 149.915 18.485 ;
        RECT 154.010 18.245 156.000 18.565 ;
        RECT 141.345 17.515 143.365 17.795 ;
        RECT 148.910 17.670 150.710 17.860 ;
        RECT 148.910 17.605 149.170 17.670 ;
        RECT 141.205 16.955 141.435 17.365 ;
        RECT 140.545 16.755 141.435 16.955 ;
        RECT 141.205 16.365 141.435 16.755 ;
        RECT 141.645 16.865 141.875 17.365 ;
        RECT 142.115 16.865 142.435 16.915 ;
        RECT 141.645 16.705 142.435 16.865 ;
        RECT 141.645 16.365 141.875 16.705 ;
        RECT 142.115 16.655 142.435 16.705 ;
        RECT 141.395 16.195 141.685 16.205 ;
        RECT 143.075 16.195 143.365 17.515 ;
        RECT 147.665 17.075 149.885 17.275 ;
        RECT 147.665 16.825 147.865 17.075 ;
        RECT 147.665 16.735 147.875 16.825 ;
        RECT 141.365 16.155 143.375 16.195 ;
        RECT 141.365 15.915 143.395 16.155 ;
        RECT 142.115 15.405 142.435 15.455 ;
        RECT 139.055 15.095 139.570 15.275 ;
        RECT 140.235 15.245 142.435 15.405 ;
        RECT 140.235 15.095 140.395 15.245 ;
        RECT 142.115 15.195 142.435 15.245 ;
        RECT 143.115 15.275 143.395 15.915 ;
        RECT 147.675 15.475 147.875 16.735 ;
        RECT 148.910 16.495 149.170 16.815 ;
        RECT 149.685 16.705 149.885 17.075 ;
        RECT 148.925 16.225 149.155 16.495 ;
        RECT 149.315 16.475 150.315 16.705 ;
        RECT 150.520 16.515 150.710 17.670 ;
        RECT 149.315 16.035 150.315 16.265 ;
        RECT 150.475 16.225 150.710 16.515 ;
        RECT 150.520 16.200 150.710 16.225 ;
        RECT 151.000 16.775 151.650 17.245 ;
        RECT 154.010 17.205 154.230 18.245 ;
        RECT 154.930 17.735 157.190 17.995 ;
        RECT 154.760 17.205 154.990 17.575 ;
        RECT 154.000 16.985 154.990 17.205 ;
        RECT 144.480 15.275 144.660 15.285 ;
        RECT 145.885 15.275 147.875 15.475 ;
        RECT 139.055 15.045 140.405 15.095 ;
        RECT 137.850 14.855 140.405 15.045 ;
        RECT 143.115 15.035 146.100 15.275 ;
        RECT 149.745 15.265 149.935 16.035 ;
        RECT 151.000 15.775 152.480 16.775 ;
        RECT 154.760 16.575 154.990 16.985 ;
        RECT 155.200 17.200 155.430 17.575 ;
        RECT 155.870 17.200 156.190 17.225 ;
        RECT 155.200 16.990 156.190 17.200 ;
        RECT 155.200 16.575 155.430 16.990 ;
        RECT 155.870 16.965 156.190 16.990 ;
        RECT 154.950 16.405 155.240 16.415 ;
        RECT 156.930 16.405 157.190 17.735 ;
        RECT 154.870 16.145 157.210 16.405 ;
        RECT 151.000 15.475 151.650 15.775 ;
        RECT 155.870 15.470 156.190 15.495 ;
        RECT 152.015 15.265 152.725 15.280 ;
        RECT 137.850 14.795 139.570 14.855 ;
        RECT 137.850 14.765 138.270 14.795 ;
        RECT 137.850 14.585 138.150 14.765 ;
        RECT 135.930 14.285 138.150 14.585 ;
        RECT 135.785 13.315 136.015 14.110 ;
        RECT 134.570 13.105 136.015 13.315 ;
        RECT 135.785 11.610 136.015 13.105 ;
        RECT 136.225 12.115 136.455 14.110 ;
        RECT 137.365 12.135 137.685 12.145 ;
        RECT 136.925 12.115 137.685 12.135 ;
        RECT 136.225 11.895 137.685 12.115 ;
        RECT 136.225 11.875 137.175 11.895 ;
        RECT 137.365 11.885 137.685 11.895 ;
        RECT 136.225 11.610 136.455 11.875 ;
        RECT 137.850 11.405 138.150 14.285 ;
        RECT 140.235 13.145 140.395 14.855 ;
        RECT 143.115 14.535 143.395 15.035 ;
        RECT 141.375 14.295 143.395 14.535 ;
        RECT 141.235 13.145 141.465 14.100 ;
        RECT 140.235 12.985 141.465 13.145 ;
        RECT 141.235 11.600 141.465 12.985 ;
        RECT 141.675 11.995 141.905 14.100 ;
        RECT 142.575 11.995 142.895 12.020 ;
        RECT 141.675 11.785 142.895 11.995 ;
        RECT 141.675 11.600 141.905 11.785 ;
        RECT 142.575 11.760 142.895 11.785 ;
        RECT 143.115 11.425 143.395 14.295 ;
        RECT 135.890 11.105 138.150 11.405 ;
        RECT 141.425 11.185 143.395 11.425 ;
        RECT 141.425 11.165 141.715 11.185 ;
        RECT 135.215 10.445 136.945 10.845 ;
        RECT 140.585 10.460 142.325 10.925 ;
        RECT 142.575 10.460 142.895 10.485 ;
        RECT 135.215 10.185 137.215 10.445 ;
        RECT 140.585 10.250 142.895 10.460 ;
        RECT 135.215 9.985 136.945 10.185 ;
        RECT 140.585 9.985 142.325 10.250 ;
        RECT 142.575 10.225 142.895 10.250 ;
        RECT 135.645 8.755 136.645 9.985 ;
        RECT 141.045 8.945 142.045 9.985 ;
        RECT 139.485 6.925 139.805 6.935 ;
        RECT 140.065 6.925 141.065 8.255 ;
        RECT 139.485 6.685 141.345 6.925 ;
        RECT 139.485 6.675 139.805 6.685 ;
        RECT 138.545 5.965 140.505 6.165 ;
        RECT 138.545 4.145 138.745 5.965 ;
        RECT 140.305 5.775 140.505 5.965 ;
        RECT 139.515 5.245 139.775 5.745 ;
        RECT 139.915 5.545 140.915 5.775 ;
        RECT 141.105 5.585 141.345 6.685 ;
        RECT 139.915 5.105 140.915 5.335 ;
        RECT 141.075 5.295 141.345 5.585 ;
        RECT 141.105 5.285 141.345 5.295 ;
        RECT 141.605 5.885 142.345 6.225 ;
        RECT 140.425 4.215 140.605 5.105 ;
        RECT 141.605 4.885 143.135 5.885 ;
        RECT 141.605 4.635 142.345 4.885 ;
        RECT 144.480 4.215 144.660 15.035 ;
        RECT 145.885 12.375 146.085 15.035 ;
        RECT 149.740 15.010 152.725 15.265 ;
        RECT 153.505 15.260 156.190 15.470 ;
        RECT 153.505 15.045 153.715 15.260 ;
        RECT 155.870 15.235 156.190 15.260 ;
        RECT 149.740 15.000 152.190 15.010 ;
        RECT 147.290 13.995 147.810 14.375 ;
        RECT 146.500 12.975 147.810 13.995 ;
        RECT 149.745 13.845 149.935 15.000 ;
        RECT 147.290 12.805 147.810 12.975 ;
        RECT 147.465 12.375 147.725 12.435 ;
        RECT 145.885 12.175 147.725 12.375 ;
        RECT 147.465 12.115 147.725 12.175 ;
        RECT 148.075 11.925 148.335 13.695 ;
        RECT 148.510 13.615 151.010 13.845 ;
        RECT 151.245 13.655 151.505 13.715 ;
        RECT 148.510 13.175 151.010 13.405 ;
        RECT 151.215 13.365 151.505 13.655 ;
        RECT 148.845 13.025 149.045 13.175 ;
        RECT 148.815 12.705 149.075 13.025 ;
        RECT 151.245 11.925 151.505 13.365 ;
        RECT 148.065 11.625 151.545 11.925 ;
        RECT 148.075 11.605 148.335 11.625 ;
        RECT 149.765 11.005 150.015 11.625 ;
        RECT 149.345 9.975 150.345 11.005 ;
        RECT 138.495 3.995 138.765 4.145 ;
        RECT 136.605 3.805 138.765 3.995 ;
        RECT 140.425 4.035 144.660 4.215 ;
        RECT 136.605 3.795 138.555 3.805 ;
        RECT 136.605 2.745 136.805 3.795 ;
        RECT 137.865 3.065 138.455 3.205 ;
        RECT 133.890 2.485 136.820 2.745 ;
        RECT 118.385 1.100 121.880 1.390 ;
        RECT 136.605 1.375 136.805 2.485 ;
        RECT 136.975 2.065 138.455 3.065 ;
        RECT 140.425 2.935 140.605 4.035 ;
        RECT 152.455 3.350 152.725 15.010 ;
        RECT 152.935 14.755 153.720 15.045 ;
        RECT 153.505 12.865 153.715 14.755 ;
        RECT 156.950 14.625 157.210 16.145 ;
        RECT 157.520 14.660 158.520 14.895 ;
        RECT 180.340 14.660 180.600 27.330 ;
        RECT 157.520 14.625 180.600 14.660 ;
        RECT 156.930 14.400 180.600 14.625 ;
        RECT 156.930 14.385 158.520 14.400 ;
        RECT 154.880 14.335 158.520 14.385 ;
        RECT 154.880 14.125 157.210 14.335 ;
        RECT 154.930 14.105 155.220 14.125 ;
        RECT 154.740 12.865 154.970 13.900 ;
        RECT 153.460 12.655 154.970 12.865 ;
        RECT 154.740 11.400 154.970 12.655 ;
        RECT 155.180 11.755 155.410 13.900 ;
        RECT 156.300 11.755 156.620 11.770 ;
        RECT 155.180 11.525 156.620 11.755 ;
        RECT 155.180 11.400 155.410 11.525 ;
        RECT 156.300 11.510 156.620 11.525 ;
        RECT 156.950 11.235 157.210 14.125 ;
        RECT 157.520 13.865 158.520 14.335 ;
        RECT 154.880 10.975 157.210 11.235 ;
        RECT 154.930 10.965 155.220 10.975 ;
        RECT 154.210 10.210 156.020 10.665 ;
        RECT 156.300 10.210 156.620 10.225 ;
        RECT 154.210 9.980 156.620 10.210 ;
        RECT 154.210 9.795 156.020 9.980 ;
        RECT 156.300 9.965 156.620 9.980 ;
        RECT 154.620 8.445 155.620 9.795 ;
        RECT 154.870 7.595 155.200 8.445 ;
        RECT 160.335 7.595 160.665 13.275 ;
        RECT 154.870 7.265 160.665 7.595 ;
        RECT 154.870 7.230 155.200 7.265 ;
        RECT 143.405 3.080 152.725 3.350 ;
        RECT 138.715 2.365 139.045 2.795 ;
        RECT 139.200 2.705 141.700 2.935 ;
        RECT 141.935 2.745 142.135 2.755 ;
        RECT 138.750 2.065 139.010 2.365 ;
        RECT 139.200 2.265 141.700 2.495 ;
        RECT 141.905 2.455 142.135 2.745 ;
        RECT 137.865 1.755 138.455 2.065 ;
        RECT 139.725 1.375 139.925 2.265 ;
        RECT 136.605 1.175 139.925 1.375 ;
        RECT 119.975 0.675 120.295 1.100 ;
        RECT 138.750 0.825 139.010 0.885 ;
        RECT 140.375 0.825 140.685 0.835 ;
        RECT 141.935 0.825 142.135 2.455 ;
        RECT 119.585 -0.355 120.585 0.675 ;
        RECT 138.750 0.625 142.135 0.825 ;
        RECT 138.750 0.565 139.010 0.625 ;
        RECT 140.375 0.195 140.685 0.625 ;
        RECT 113.605 -3.450 140.550 -3.380 ;
        RECT 143.405 -3.450 143.675 3.080 ;
        RECT 113.605 -3.650 143.675 -3.450 ;
        RECT 140.175 -3.720 143.675 -3.650 ;
        RECT 6.830 -5.190 38.280 -4.780 ;
        RECT 35.320 -5.220 38.280 -5.190 ;
      LAYER met2 ;
        RECT 72.900 87.700 73.420 87.730 ;
        RECT 72.900 87.180 77.705 87.700 ;
        RECT 72.900 87.150 73.420 87.180 ;
        RECT 72.320 72.900 73.320 72.930 ;
        RECT 72.320 71.900 78.840 72.900 ;
        RECT 72.320 71.870 73.320 71.900 ;
        RECT 59.425 63.910 59.895 63.930 ;
        RECT 59.400 63.390 62.100 63.910 ;
        RECT 59.425 63.370 59.895 63.390 ;
        RECT 68.640 62.420 69.160 66.790 ;
        RECT 68.610 61.900 69.190 62.420 ;
        RECT 64.290 47.480 64.810 47.510 ;
        RECT 62.365 46.960 64.810 47.480 ;
        RECT 64.290 46.930 64.810 46.960 ;
        RECT 138.345 44.515 138.675 44.545 ;
        RECT 138.345 44.185 160.665 44.515 ;
        RECT 138.345 44.155 138.675 44.185 ;
        RECT 104.620 43.610 104.940 43.870 ;
        RECT 104.680 42.370 104.880 43.610 ;
        RECT 104.620 42.110 104.940 42.370 ;
        RECT 124.955 41.535 125.245 43.395 ;
        RECT 153.555 43.240 153.875 43.500 ;
        RECT 153.615 42.000 153.815 43.240 ;
        RECT 153.555 41.740 153.875 42.000 ;
        RECT 124.925 41.245 125.275 41.535 ;
        RECT 103.855 38.750 104.175 39.010 ;
        RECT 103.885 37.500 104.145 38.750 ;
        RECT 152.790 38.380 153.110 38.640 ;
        RECT 124.055 37.860 124.395 38.140 ;
        RECT 124.085 36.800 124.365 37.860 ;
        RECT 152.820 37.130 153.080 38.380 ;
        RECT 87.070 34.210 87.330 34.530 ;
        RECT 119.380 34.335 119.640 34.655 ;
        RECT 106.475 34.270 106.735 34.310 ;
        RECT 87.085 32.985 87.315 34.210 ;
        RECT 100.795 33.950 101.055 34.270 ;
        RECT 106.015 34.030 106.735 34.270 ;
        RECT 87.070 32.665 87.330 32.985 ;
        RECT 100.820 32.735 101.030 33.950 ;
        RECT 100.795 32.415 101.055 32.735 ;
        RECT 106.015 32.610 106.255 34.030 ;
        RECT 106.475 33.990 106.735 34.030 ;
        RECT 12.080 32.130 12.400 32.390 ;
        RECT 95.905 32.290 96.225 32.320 ;
        RECT 106.005 32.290 106.265 32.610 ;
        RECT 12.110 31.020 12.370 32.130 ;
        RECT 94.615 32.090 96.225 32.290 ;
        RECT 94.615 31.730 94.815 32.090 ;
        RECT 95.905 32.060 96.225 32.090 ;
        RECT 115.025 31.820 115.325 33.450 ;
        RECT 119.415 32.510 119.605 34.335 ;
        RECT 119.350 32.250 119.670 32.510 ;
        RECT 124.255 32.320 124.515 34.590 ;
        RECT 136.005 33.840 136.265 34.160 ;
        RECT 155.410 33.900 155.670 33.940 ;
        RECT 136.020 32.615 136.250 33.840 ;
        RECT 149.730 33.580 149.990 33.900 ;
        RECT 154.950 33.660 155.670 33.900 ;
        RECT 136.005 32.295 136.265 32.615 ;
        RECT 149.755 32.365 149.965 33.580 ;
        RECT 149.730 32.045 149.990 32.365 ;
        RECT 154.950 32.240 155.190 33.660 ;
        RECT 155.410 33.620 155.670 33.660 ;
        RECT 144.840 31.920 145.160 31.950 ;
        RECT 154.940 31.920 155.200 32.240 ;
        RECT 94.555 31.470 94.875 31.730 ;
        RECT 114.995 31.520 115.355 31.820 ;
        RECT 143.550 31.720 145.160 31.920 ;
        RECT 143.550 31.360 143.750 31.720 ;
        RECT 144.840 31.690 145.160 31.720 ;
        RECT 13.380 31.310 13.640 31.340 ;
        RECT 13.380 31.050 14.950 31.310 ;
        RECT 143.490 31.100 143.810 31.360 ;
        RECT 13.380 31.020 13.640 31.050 ;
        RECT 13.820 29.300 14.080 29.620 ;
        RECT 119.785 29.370 120.045 29.690 ;
        RECT 13.870 28.010 14.030 29.300 ;
        RECT 87.500 28.940 87.760 29.260 ;
        RECT 101.255 28.980 101.515 29.300 ;
        RECT 13.790 27.750 14.110 28.010 ;
        RECT 23.650 27.680 23.970 27.940 ;
        RECT 25.670 27.890 25.990 28.150 ;
        RECT 23.695 26.030 23.925 27.680 ;
        RECT 25.740 26.920 25.920 27.890 ;
        RECT 87.525 27.530 87.735 28.940 ;
        RECT 94.460 27.680 94.780 27.940 ;
        RECT 101.305 27.840 101.465 28.980 ;
        RECT 106.720 28.810 106.980 29.130 ;
        RECT 87.500 27.210 87.760 27.530 ;
        RECT 25.700 26.600 25.960 26.920 ;
        RECT 94.525 26.830 94.715 27.680 ;
        RECT 101.255 27.520 101.515 27.840 ;
        RECT 106.745 27.450 106.955 28.810 ;
        RECT 114.275 28.240 114.595 28.500 ;
        RECT 114.315 27.590 114.555 28.240 ;
        RECT 119.790 27.970 120.040 29.370 ;
        RECT 119.755 27.710 120.075 27.970 ;
        RECT 106.720 27.130 106.980 27.450 ;
        RECT 114.305 27.270 114.565 27.590 ;
        RECT 124.925 27.390 125.185 29.450 ;
        RECT 136.435 28.570 136.695 28.890 ;
        RECT 150.190 28.610 150.450 28.930 ;
        RECT 136.460 27.160 136.670 28.570 ;
        RECT 143.395 27.310 143.715 27.570 ;
        RECT 150.240 27.470 150.400 28.610 ;
        RECT 155.655 28.440 155.915 28.760 ;
        RECT 136.435 26.840 136.695 27.160 ;
        RECT 94.460 26.570 94.780 26.830 ;
        RECT 143.460 26.460 143.650 27.310 ;
        RECT 150.190 27.150 150.450 27.470 ;
        RECT 155.680 27.080 155.890 28.440 ;
        RECT 155.655 26.760 155.915 27.080 ;
        RECT 143.395 26.200 143.715 26.460 ;
        RECT 23.650 25.770 23.970 26.030 ;
        RECT 11.250 25.590 11.510 25.670 ;
        RECT 12.410 25.590 12.730 25.640 ;
        RECT 1.130 25.230 1.390 25.550 ;
        RECT 11.250 25.430 12.730 25.590 ;
        RECT 11.250 25.350 11.510 25.430 ;
        RECT 12.410 25.380 12.730 25.430 ;
        RECT 1.150 24.160 1.370 25.230 ;
        RECT 1.130 23.840 1.390 24.160 ;
        RECT 8.820 22.000 9.100 22.030 ;
        RECT 7.670 21.720 9.100 22.000 ;
        RECT 8.820 21.690 9.100 21.720 ;
        RECT 14.860 18.780 15.180 19.040 ;
        RECT 14.920 17.370 15.120 18.780 ;
        RECT 148.880 17.635 149.200 17.895 ;
        RECT 14.890 17.050 15.150 17.370 ;
        RECT 118.475 15.015 118.735 17.075 ;
        RECT 129.095 16.875 129.355 17.195 ;
        RECT 136.680 17.015 136.940 17.335 ;
        RECT 123.585 16.495 123.905 16.755 ;
        RECT 123.620 15.095 123.870 16.495 ;
        RECT 129.105 16.225 129.345 16.875 ;
        RECT 129.065 15.965 129.385 16.225 ;
        RECT 136.705 15.655 136.915 17.015 ;
        RECT 142.145 16.625 142.405 16.945 ;
        RECT 148.945 16.785 149.135 17.635 ;
        RECT 155.900 16.935 156.160 17.255 ;
        RECT 136.680 15.335 136.940 15.655 ;
        RECT 142.195 15.485 142.355 16.625 ;
        RECT 148.880 16.525 149.200 16.785 ;
        RECT 155.925 15.525 156.135 16.935 ;
        RECT 142.145 15.165 142.405 15.485 ;
        RECT 155.900 15.205 156.160 15.525 ;
        RECT 123.615 14.775 123.875 15.095 ;
        RECT 160.335 13.245 160.665 44.185 ;
        RECT 173.890 41.165 174.180 43.025 ;
        RECT 173.860 40.875 174.210 41.165 ;
        RECT 172.990 37.490 173.330 37.770 ;
        RECT 173.020 36.430 173.300 37.490 ;
        RECT 168.315 33.965 168.575 34.285 ;
        RECT 163.960 31.450 164.260 33.080 ;
        RECT 168.350 32.140 168.540 33.965 ;
        RECT 168.285 31.880 168.605 32.140 ;
        RECT 173.190 31.950 173.450 34.220 ;
        RECT 163.930 31.150 164.290 31.450 ;
        RECT 168.720 29.000 168.980 29.320 ;
        RECT 163.210 27.870 163.530 28.130 ;
        RECT 163.250 27.220 163.490 27.870 ;
        RECT 168.725 27.600 168.975 29.000 ;
        RECT 168.690 27.340 169.010 27.600 ;
        RECT 163.240 26.900 163.500 27.220 ;
        RECT 173.860 27.020 174.120 29.080 ;
        RECT 128.305 12.645 128.665 12.945 ;
        RECT 148.785 12.735 149.105 12.995 ;
        RECT 160.305 12.915 160.695 13.245 ;
        RECT 17.060 12.020 17.380 12.280 ;
        RECT 12.330 11.810 12.590 11.880 ;
        RECT 13.250 11.810 13.570 11.850 ;
        RECT 12.330 11.630 13.570 11.810 ;
        RECT 12.330 11.560 12.590 11.630 ;
        RECT 13.250 11.590 13.570 11.630 ;
        RECT 17.130 11.250 17.310 12.020 ;
        RECT 50.320 11.890 50.580 11.935 ;
        RECT 52.690 11.890 53.010 11.905 ;
        RECT 50.320 11.660 53.010 11.890 ;
        RECT 50.320 11.615 50.580 11.660 ;
        RECT 52.690 11.645 53.010 11.660 ;
        RECT 58.880 11.890 59.140 11.935 ;
        RECT 60.380 11.890 60.700 11.905 ;
        RECT 58.880 11.660 60.700 11.890 ;
        RECT 58.880 11.615 59.140 11.660 ;
        RECT 60.380 11.645 60.700 11.660 ;
        RECT 66.700 11.890 66.960 11.935 ;
        RECT 67.820 11.890 68.140 11.905 ;
        RECT 66.700 11.660 68.140 11.890 ;
        RECT 66.700 11.615 66.960 11.660 ;
        RECT 67.820 11.645 68.140 11.660 ;
        RECT 74.620 11.890 74.940 11.905 ;
        RECT 75.740 11.890 76.060 11.905 ;
        RECT 74.620 11.660 76.060 11.890 ;
        RECT 74.620 11.645 74.940 11.660 ;
        RECT 75.740 11.645 76.060 11.660 ;
        RECT 82.290 11.890 82.550 11.935 ;
        RECT 83.610 11.890 83.930 11.905 ;
        RECT 82.290 11.660 83.930 11.890 ;
        RECT 82.290 11.615 82.550 11.660 ;
        RECT 83.610 11.645 83.930 11.660 ;
        RECT 90.220 11.890 90.480 11.935 ;
        RECT 91.370 11.890 91.690 11.905 ;
        RECT 90.220 11.660 91.690 11.890 ;
        RECT 90.220 11.615 90.480 11.660 ;
        RECT 91.370 11.645 91.690 11.660 ;
        RECT 97.450 11.890 97.710 11.935 ;
        RECT 98.470 11.890 98.790 11.905 ;
        RECT 97.450 11.660 98.790 11.890 ;
        RECT 97.450 11.615 97.710 11.660 ;
        RECT 98.470 11.645 98.790 11.660 ;
        RECT 17.090 10.930 17.350 11.250 ;
        RECT 1.870 10.640 2.190 10.900 ;
        RECT 53.700 10.845 53.960 11.165 ;
        RECT 61.290 10.895 61.550 11.215 ;
        RECT 68.900 10.915 69.160 11.235 ;
        RECT 1.935 9.870 2.125 10.640 ;
        RECT 12.200 10.390 12.520 10.650 ;
        RECT 1.900 9.550 2.160 9.870 ;
        RECT 12.270 9.710 12.450 10.390 ;
        RECT 12.230 9.390 12.490 9.710 ;
        RECT 53.710 9.625 53.950 10.845 ;
        RECT 53.710 9.375 54.260 9.625 ;
        RECT 55.650 9.530 55.910 9.850 ;
        RECT 61.300 9.675 61.540 10.895 ;
        RECT 53.940 9.365 54.260 9.375 ;
        RECT 55.695 8.315 55.865 9.530 ;
        RECT 61.300 9.425 61.850 9.675 ;
        RECT 63.240 9.580 63.500 9.900 ;
        RECT 68.910 9.695 69.150 10.915 ;
        RECT 76.900 10.875 77.160 11.195 ;
        RECT 84.710 10.895 84.970 11.215 ;
        RECT 61.530 9.415 61.850 9.425 ;
        RECT 63.285 8.365 63.455 9.580 ;
        RECT 68.910 9.445 69.460 9.695 ;
        RECT 70.850 9.600 71.110 9.920 ;
        RECT 76.910 9.655 77.150 10.875 ;
        RECT 69.140 9.435 69.460 9.445 ;
        RECT 70.895 8.385 71.065 9.600 ;
        RECT 76.910 9.405 77.460 9.655 ;
        RECT 78.850 9.560 79.110 9.880 ;
        RECT 84.720 9.675 84.960 10.895 ;
        RECT 92.300 10.875 92.560 11.195 ;
        RECT 77.140 9.395 77.460 9.405 ;
        RECT 54.350 8.175 55.865 8.315 ;
        RECT 9.020 7.400 9.340 7.405 ;
        RECT 10.130 7.400 10.390 7.435 ;
        RECT 9.020 7.150 10.390 7.400 ;
        RECT 9.020 7.145 9.340 7.150 ;
        RECT 10.130 7.115 10.390 7.150 ;
        RECT 54.350 6.825 54.490 8.175 ;
        RECT 55.695 8.160 55.865 8.175 ;
        RECT 61.940 8.225 63.455 8.365 ;
        RECT 61.940 6.875 62.080 8.225 ;
        RECT 63.285 8.210 63.455 8.225 ;
        RECT 69.550 8.245 71.065 8.385 ;
        RECT 78.895 8.345 79.065 9.560 ;
        RECT 84.720 9.425 85.270 9.675 ;
        RECT 86.660 9.580 86.920 9.900 ;
        RECT 92.310 9.655 92.550 10.875 ;
        RECT 99.690 10.845 99.950 11.165 ;
        RECT 84.950 9.415 85.270 9.425 ;
        RECT 86.705 8.365 86.875 9.580 ;
        RECT 92.310 9.405 92.860 9.655 ;
        RECT 94.250 9.560 94.510 9.880 ;
        RECT 99.700 9.625 99.940 10.845 ;
        RECT 119.145 9.875 119.405 12.145 ;
        RECT 123.990 11.955 124.310 12.215 ;
        RECT 124.055 10.130 124.245 11.955 ;
        RECT 128.335 11.015 128.635 12.645 ;
        RECT 147.435 12.375 147.755 12.405 ;
        RECT 148.845 12.375 149.045 12.735 ;
        RECT 147.435 12.175 149.045 12.375 ;
        RECT 137.395 11.855 137.655 12.175 ;
        RECT 147.435 12.145 147.755 12.175 ;
        RECT 136.925 10.435 137.185 10.475 ;
        RECT 137.405 10.435 137.645 11.855 ;
        RECT 142.605 11.730 142.865 12.050 ;
        RECT 142.630 10.515 142.840 11.730 ;
        RECT 156.330 11.480 156.590 11.800 ;
        RECT 136.925 10.195 137.645 10.435 ;
        RECT 142.605 10.195 142.865 10.515 ;
        RECT 156.345 10.255 156.575 11.480 ;
        RECT 136.925 10.155 137.185 10.195 ;
        RECT 92.540 9.395 92.860 9.405 ;
        RECT 69.550 6.895 69.690 8.245 ;
        RECT 70.895 8.230 71.065 8.245 ;
        RECT 77.550 8.205 79.065 8.345 ;
        RECT 54.290 6.505 54.550 6.825 ;
        RECT 61.880 6.555 62.140 6.875 ;
        RECT 69.490 6.575 69.750 6.895 ;
        RECT 77.550 6.855 77.690 8.205 ;
        RECT 78.895 8.190 79.065 8.205 ;
        RECT 85.360 8.225 86.875 8.365 ;
        RECT 94.295 8.345 94.465 9.560 ;
        RECT 99.700 9.375 100.250 9.625 ;
        RECT 101.640 9.530 101.900 9.850 ;
        RECT 124.020 9.810 124.280 10.130 ;
        RECT 156.330 9.935 156.590 10.255 ;
        RECT 99.930 9.365 100.250 9.375 ;
        RECT 85.360 6.875 85.500 8.225 ;
        RECT 86.705 8.210 86.875 8.225 ;
        RECT 92.950 8.205 94.465 8.345 ;
        RECT 101.685 8.315 101.855 9.530 ;
        RECT 106.230 8.685 106.490 9.005 ;
        RECT 77.490 6.535 77.750 6.855 ;
        RECT 85.300 6.555 85.560 6.875 ;
        RECT 92.950 6.855 93.090 8.205 ;
        RECT 94.295 8.190 94.465 8.205 ;
        RECT 100.340 8.175 101.855 8.315 ;
        RECT 92.890 6.535 93.150 6.855 ;
        RECT 100.340 6.825 100.480 8.175 ;
        RECT 101.685 8.160 101.855 8.175 ;
        RECT 106.270 7.495 106.450 8.685 ;
        RECT 106.200 7.235 106.520 7.495 ;
        RECT 100.280 6.505 100.540 6.825 ;
        RECT 119.295 6.605 119.575 7.665 ;
        RECT 119.265 6.325 119.605 6.605 ;
        RECT 139.515 5.715 139.775 6.965 ;
        RECT 139.485 5.455 139.805 5.715 ;
        RECT 17.090 5.090 17.350 5.410 ;
        RECT 106.430 5.135 106.690 5.455 ;
        RECT 17.130 4.130 17.310 5.090 ;
        RECT 54.000 4.575 54.260 4.895 ;
        RECT 61.590 4.625 61.850 4.945 ;
        RECT 69.200 4.645 69.460 4.965 ;
        RECT 17.090 3.810 17.350 4.130 ;
        RECT 45.340 4.125 45.600 4.445 ;
        RECT 45.365 3.235 45.575 4.125 ;
        RECT 54.040 3.875 54.220 4.575 ;
        RECT 61.630 3.925 61.810 4.625 ;
        RECT 69.240 3.945 69.420 4.645 ;
        RECT 77.200 4.605 77.460 4.925 ;
        RECT 85.010 4.625 85.270 4.945 ;
        RECT 53.970 3.615 54.290 3.875 ;
        RECT 61.560 3.665 61.880 3.925 ;
        RECT 69.170 3.685 69.490 3.945 ;
        RECT 77.240 3.905 77.420 4.605 ;
        RECT 85.050 3.925 85.230 4.625 ;
        RECT 92.600 4.605 92.860 4.925 ;
        RECT 77.170 3.645 77.490 3.905 ;
        RECT 84.980 3.665 85.300 3.925 ;
        RECT 92.640 3.905 92.820 4.605 ;
        RECT 99.990 4.575 100.250 4.895 ;
        RECT 92.570 3.645 92.890 3.905 ;
        RECT 100.030 3.875 100.210 4.575 ;
        RECT 106.465 4.225 106.655 5.135 ;
        RECT 106.400 3.965 106.720 4.225 ;
        RECT 99.960 3.615 100.280 3.875 ;
        RECT 45.340 2.915 45.600 3.235 ;
        RECT 118.385 2.930 118.735 3.220 ;
        RECT 25.975 2.160 26.295 2.420 ;
        RECT 26.040 1.250 26.230 2.160 ;
        RECT 54.100 1.945 54.360 2.265 ;
        RECT 61.690 1.995 61.950 2.315 ;
        RECT 69.300 2.015 69.560 2.335 ;
        RECT 54.145 1.425 54.315 1.945 ;
        RECT 61.735 1.475 61.905 1.995 ;
        RECT 69.345 1.495 69.515 2.015 ;
        RECT 77.300 1.975 77.560 2.295 ;
        RECT 85.110 1.995 85.370 2.315 ;
        RECT 26.005 0.930 26.265 1.250 ;
        RECT 54.100 1.105 54.360 1.425 ;
        RECT 61.690 1.155 61.950 1.475 ;
        RECT 69.300 1.175 69.560 1.495 ;
        RECT 77.345 1.455 77.515 1.975 ;
        RECT 85.155 1.475 85.325 1.995 ;
        RECT 92.700 1.975 92.960 2.295 ;
        RECT 77.300 1.135 77.560 1.455 ;
        RECT 85.110 1.155 85.370 1.475 ;
        RECT 92.745 1.455 92.915 1.975 ;
        RECT 100.090 1.945 100.350 2.265 ;
        RECT 92.700 1.135 92.960 1.455 ;
        RECT 100.135 1.425 100.305 1.945 ;
        RECT 100.090 1.105 100.350 1.425 ;
        RECT 118.415 1.070 118.705 2.930 ;
        RECT 138.720 2.095 139.040 2.355 ;
        RECT 138.780 0.855 138.980 2.095 ;
        RECT 138.720 0.595 139.040 0.855 ;
        RECT 48.970 -0.385 49.230 -0.345 ;
        RECT 50.160 -0.385 50.480 -0.375 ;
        RECT 48.970 -0.625 50.480 -0.385 ;
        RECT 48.970 -0.665 49.230 -0.625 ;
        RECT 50.160 -0.635 50.480 -0.625 ;
        RECT 51.830 -0.385 52.090 -0.345 ;
        RECT 52.930 -0.385 53.250 -0.375 ;
        RECT 51.830 -0.625 53.250 -0.385 ;
        RECT 51.830 -0.665 52.090 -0.625 ;
        RECT 52.930 -0.635 53.250 -0.625 ;
        RECT 59.400 -0.385 59.660 -0.345 ;
        RECT 60.530 -0.385 60.850 -0.375 ;
        RECT 59.400 -0.625 60.850 -0.385 ;
        RECT 59.400 -0.665 59.660 -0.625 ;
        RECT 60.530 -0.635 60.850 -0.625 ;
        RECT 67.010 -0.385 67.270 -0.345 ;
        RECT 68.330 -0.385 68.650 -0.375 ;
        RECT 67.010 -0.625 68.650 -0.385 ;
        RECT 67.010 -0.665 67.270 -0.625 ;
        RECT 68.330 -0.635 68.650 -0.625 ;
        RECT 74.890 -0.385 75.150 -0.345 ;
        RECT 76.310 -0.385 76.630 -0.375 ;
        RECT 74.890 -0.625 76.630 -0.385 ;
        RECT 74.890 -0.665 75.150 -0.625 ;
        RECT 76.310 -0.635 76.630 -0.625 ;
        RECT 82.760 -0.385 83.020 -0.345 ;
        RECT 83.970 -0.385 84.290 -0.375 ;
        RECT 82.760 -0.625 84.290 -0.385 ;
        RECT 82.760 -0.665 83.020 -0.625 ;
        RECT 83.970 -0.635 84.290 -0.625 ;
        RECT 90.700 -0.385 90.960 -0.345 ;
        RECT 91.840 -0.385 92.160 -0.375 ;
        RECT 90.700 -0.625 92.160 -0.385 ;
        RECT 90.700 -0.665 90.960 -0.625 ;
        RECT 91.840 -0.635 92.160 -0.625 ;
        RECT 97.950 -0.385 98.210 -0.345 ;
        RECT 99.110 -0.385 99.430 -0.375 ;
        RECT 97.950 -0.625 99.430 -0.385 ;
        RECT 97.950 -0.665 98.210 -0.625 ;
        RECT 99.110 -0.635 99.430 -0.625 ;
        RECT 103.570 -0.385 103.830 -0.345 ;
        RECT 105.630 -0.385 105.950 -0.375 ;
        RECT 103.570 -0.625 105.950 -0.385 ;
        RECT 103.570 -0.665 103.830 -0.625 ;
        RECT 105.630 -0.635 105.950 -0.625 ;
        RECT 50.675 -1.595 50.945 -1.565 ;
        RECT 47.985 -1.865 50.945 -1.595 ;
        RECT 50.675 -1.895 50.945 -1.865 ;
      LAYER met3 ;
        RECT -322.220 410.650 -291.820 442.510 ;
        RECT -290.620 410.650 -260.220 442.510 ;
        RECT -259.020 410.650 -228.620 442.510 ;
        RECT -227.420 410.650 -197.020 442.510 ;
        RECT -195.820 410.650 -165.420 442.510 ;
        RECT -164.220 410.650 -133.820 442.510 ;
        RECT -132.620 410.650 -102.220 442.510 ;
        RECT -101.020 410.650 -70.620 442.510 ;
        RECT -69.420 410.650 -39.020 442.510 ;
        RECT -37.820 410.650 -7.420 442.510 ;
        RECT -6.220 410.650 24.180 442.510 ;
        RECT 25.380 410.650 55.780 442.510 ;
        RECT -324.780 392.785 -324.260 395.750 ;
        RECT -324.805 392.275 -324.235 392.785 ;
        RECT -324.780 392.270 -324.260 392.275 ;
        RECT -322.220 377.590 -291.820 409.450 ;
        RECT -290.620 377.590 -260.220 409.450 ;
        RECT -259.020 377.590 -228.620 409.450 ;
        RECT -227.420 377.590 -197.020 409.450 ;
        RECT -195.820 377.590 -165.420 409.450 ;
        RECT -164.220 377.590 -133.820 409.450 ;
        RECT -132.620 377.590 -102.220 409.450 ;
        RECT -101.020 377.590 -70.620 409.450 ;
        RECT -69.420 377.590 -39.020 409.450 ;
        RECT -37.820 377.590 -7.420 409.450 ;
        RECT -6.220 377.590 24.180 409.450 ;
        RECT 25.380 377.590 55.780 409.450 ;
        RECT -322.220 344.530 -291.820 376.390 ;
        RECT -290.620 344.530 -260.220 376.390 ;
        RECT -259.020 344.530 -228.620 376.390 ;
        RECT -227.420 344.530 -197.020 376.390 ;
        RECT -195.820 344.530 -165.420 376.390 ;
        RECT -164.220 344.530 -133.820 376.390 ;
        RECT -132.620 344.530 -102.220 376.390 ;
        RECT -101.020 344.530 -70.620 376.390 ;
        RECT -69.420 344.530 -39.020 376.390 ;
        RECT -37.820 344.530 -7.420 376.390 ;
        RECT -6.220 344.530 24.180 376.390 ;
        RECT 25.380 344.530 55.780 376.390 ;
        RECT 56.800 359.210 57.320 362.780 ;
        RECT 56.805 359.185 57.315 359.210 ;
        RECT -323.910 327.005 -323.390 329.280 ;
        RECT -323.935 326.495 -323.365 327.005 ;
        RECT -323.910 326.490 -323.390 326.495 ;
        RECT -322.220 311.470 -291.820 343.330 ;
        RECT -290.620 311.470 -260.220 343.330 ;
        RECT -259.020 311.470 -228.620 343.330 ;
        RECT -227.420 311.470 -197.020 343.330 ;
        RECT -195.820 311.470 -165.420 343.330 ;
        RECT -164.220 311.470 -133.820 343.330 ;
        RECT -132.620 311.470 -102.220 343.330 ;
        RECT -101.020 311.470 -70.620 343.330 ;
        RECT -69.420 311.470 -39.020 343.330 ;
        RECT -37.820 311.470 -7.420 343.330 ;
        RECT -6.220 311.470 24.180 343.330 ;
        RECT 25.380 311.470 55.780 343.330 ;
        RECT -322.220 278.410 -291.820 310.270 ;
        RECT -290.620 278.410 -260.220 310.270 ;
        RECT -259.020 278.410 -228.620 310.270 ;
        RECT -227.420 278.410 -197.020 310.270 ;
        RECT -195.820 278.410 -165.420 310.270 ;
        RECT -164.220 278.410 -133.820 310.270 ;
        RECT -132.620 278.410 -102.220 310.270 ;
        RECT -101.020 278.410 -70.620 310.270 ;
        RECT -69.420 278.410 -39.020 310.270 ;
        RECT -37.820 278.410 -7.420 310.270 ;
        RECT -6.220 278.410 24.180 310.270 ;
        RECT 25.380 278.410 55.780 310.270 ;
        RECT 56.850 293.925 57.370 297.260 ;
        RECT 56.825 293.415 57.395 293.925 ;
        RECT 56.850 293.410 57.370 293.415 ;
        RECT -324.060 260.875 -323.540 263.300 ;
        RECT -324.085 260.365 -323.515 260.875 ;
        RECT -324.060 260.360 -323.540 260.365 ;
        RECT -322.220 245.350 -291.820 277.210 ;
        RECT -290.620 245.350 -260.220 277.210 ;
        RECT -259.020 245.350 -228.620 277.210 ;
        RECT -227.420 245.350 -197.020 277.210 ;
        RECT -195.820 245.350 -165.420 277.210 ;
        RECT -164.220 245.350 -133.820 277.210 ;
        RECT -132.620 245.350 -102.220 277.210 ;
        RECT -101.020 245.350 -70.620 277.210 ;
        RECT -69.420 245.350 -39.020 277.210 ;
        RECT -37.820 245.350 -7.420 277.210 ;
        RECT -6.220 245.350 24.180 277.210 ;
        RECT 25.380 245.350 55.780 277.210 ;
        RECT -322.220 212.290 -291.820 244.150 ;
        RECT -290.620 212.290 -260.220 244.150 ;
        RECT -259.020 212.290 -228.620 244.150 ;
        RECT -227.420 212.290 -197.020 244.150 ;
        RECT -195.820 212.290 -165.420 244.150 ;
        RECT -164.220 212.290 -133.820 244.150 ;
        RECT -132.620 212.290 -102.220 244.150 ;
        RECT -101.020 212.290 -70.620 244.150 ;
        RECT -69.420 212.290 -39.020 244.150 ;
        RECT -37.820 212.290 -7.420 244.150 ;
        RECT -6.220 212.290 24.180 244.150 ;
        RECT 25.380 212.290 55.780 244.150 ;
        RECT 56.890 227.685 57.410 230.450 ;
        RECT 56.865 227.175 57.435 227.685 ;
        RECT 56.890 227.170 57.410 227.175 ;
        RECT 92.755 214.320 96.625 214.325 ;
        RECT 92.730 213.795 96.625 214.320 ;
        RECT 97.830 213.800 128.230 245.660 ;
        RECT 129.430 213.800 159.830 245.660 ;
        RECT 161.030 213.800 191.430 245.660 ;
        RECT 192.630 213.800 223.030 245.660 ;
        RECT 224.230 213.800 254.630 245.660 ;
        RECT 92.755 213.790 96.625 213.795 ;
        RECT -324.460 194.290 -323.940 197.380 ;
        RECT -324.455 194.265 -323.945 194.290 ;
        RECT -322.220 179.230 -291.820 211.090 ;
        RECT -290.620 179.230 -260.220 211.090 ;
        RECT -259.020 179.230 -228.620 211.090 ;
        RECT -227.420 179.230 -197.020 211.090 ;
        RECT -195.820 179.230 -165.420 211.090 ;
        RECT -164.220 179.230 -133.820 211.090 ;
        RECT -132.620 179.230 -102.220 211.090 ;
        RECT -101.020 179.230 -70.620 211.090 ;
        RECT -69.420 179.230 -39.020 211.090 ;
        RECT -37.820 179.230 -7.420 211.090 ;
        RECT -6.220 179.230 24.180 211.090 ;
        RECT 25.380 179.230 55.780 211.090 ;
        RECT 97.830 180.740 128.230 212.600 ;
        RECT 129.430 180.740 159.830 212.600 ;
        RECT 161.030 180.740 191.430 212.600 ;
        RECT 192.630 180.740 223.030 212.600 ;
        RECT 224.230 180.740 254.630 212.600 ;
        RECT -322.220 146.170 -291.820 178.030 ;
        RECT -290.620 146.170 -260.220 178.030 ;
        RECT -259.020 146.170 -228.620 178.030 ;
        RECT -227.420 146.170 -197.020 178.030 ;
        RECT -195.820 146.170 -165.420 178.030 ;
        RECT -164.220 146.170 -133.820 178.030 ;
        RECT -132.620 146.170 -102.220 178.030 ;
        RECT -101.020 146.170 -70.620 178.030 ;
        RECT -69.420 146.170 -39.020 178.030 ;
        RECT -37.820 146.170 -7.420 178.030 ;
        RECT -6.220 146.170 24.180 178.030 ;
        RECT 25.380 146.170 55.780 178.030 ;
        RECT 57.080 161.765 57.600 164.340 ;
        RECT 57.055 161.255 57.625 161.765 ;
        RECT 57.080 161.250 57.600 161.255 ;
        RECT 97.830 147.680 128.230 179.540 ;
        RECT 129.430 147.680 159.830 179.540 ;
        RECT 161.030 147.680 191.430 179.540 ;
        RECT 192.630 147.680 223.030 179.540 ;
        RECT 224.230 147.680 254.630 179.540 ;
        RECT -324.240 128.735 -323.720 131.250 ;
        RECT -324.265 128.225 -323.695 128.735 ;
        RECT -324.240 128.220 -323.720 128.225 ;
        RECT -322.220 113.110 -291.820 144.970 ;
        RECT -290.620 113.110 -260.220 144.970 ;
        RECT -259.020 113.110 -228.620 144.970 ;
        RECT -227.420 113.110 -197.020 144.970 ;
        RECT -195.820 113.110 -165.420 144.970 ;
        RECT -164.220 113.110 -133.820 144.970 ;
        RECT -132.620 113.110 -102.220 144.970 ;
        RECT -101.020 113.110 -70.620 144.970 ;
        RECT -69.420 113.110 -39.020 144.970 ;
        RECT -37.820 113.110 -7.420 144.970 ;
        RECT -6.220 113.110 24.180 144.970 ;
        RECT 25.380 113.110 55.780 144.970 ;
        RECT 95.640 129.975 96.160 133.080 ;
        RECT 95.615 129.465 96.185 129.975 ;
        RECT 95.640 129.460 96.160 129.465 ;
        RECT 97.830 114.620 128.230 146.480 ;
        RECT 129.430 114.620 159.830 146.480 ;
        RECT 161.030 114.620 191.430 146.480 ;
        RECT 192.630 114.620 223.030 146.480 ;
        RECT 224.230 114.620 254.630 146.480 ;
        RECT 255.600 115.155 258.810 115.160 ;
        RECT 255.600 114.645 258.835 115.155 ;
        RECT 255.600 114.640 258.810 114.645 ;
        RECT -322.220 80.050 -291.820 111.910 ;
        RECT -290.620 80.050 -260.220 111.910 ;
        RECT -259.020 80.050 -228.620 111.910 ;
        RECT -227.420 80.050 -197.020 111.910 ;
        RECT -195.820 80.050 -165.420 111.910 ;
        RECT -164.220 80.050 -133.820 111.910 ;
        RECT -132.620 80.050 -102.220 111.910 ;
        RECT -101.020 80.050 -70.620 111.910 ;
        RECT -69.420 80.050 -39.020 111.910 ;
        RECT -37.820 80.050 -7.420 111.910 ;
        RECT -6.220 80.050 24.180 111.910 ;
        RECT 25.380 80.050 55.780 111.910 ;
        RECT 57.120 95.695 57.640 98.050 ;
        RECT 57.095 95.185 57.665 95.695 ;
        RECT 57.120 95.180 57.640 95.185 ;
        RECT 77.115 87.700 77.685 87.725 ;
        RECT 77.115 87.180 83.470 87.700 ;
        RECT 77.115 87.155 77.685 87.180 ;
        RECT 97.830 81.560 128.230 113.420 ;
        RECT 129.430 81.560 159.830 113.420 ;
        RECT 161.030 81.560 191.430 113.420 ;
        RECT 192.630 81.560 223.030 113.420 ;
        RECT 224.230 81.560 254.630 113.420 ;
        RECT -325.110 62.395 -324.590 66.000 ;
        RECT -325.135 61.885 -324.565 62.395 ;
        RECT -325.110 61.880 -324.590 61.885 ;
        RECT -322.220 46.990 -291.820 78.850 ;
        RECT -290.620 46.990 -260.220 78.850 ;
        RECT -259.020 46.990 -228.620 78.850 ;
        RECT -227.420 46.990 -197.020 78.850 ;
        RECT -195.820 46.990 -165.420 78.850 ;
        RECT -164.220 46.990 -133.820 78.850 ;
        RECT -132.620 46.990 -102.220 78.850 ;
        RECT -101.020 46.990 -70.620 78.850 ;
        RECT -69.420 46.990 -39.020 78.850 ;
        RECT -37.820 46.990 -7.420 78.850 ;
        RECT -6.220 46.990 24.180 78.850 ;
        RECT 25.380 46.990 55.780 78.850 ;
        RECT 57.145 63.910 57.655 63.935 ;
        RECT 57.140 63.390 59.920 63.910 ;
        RECT 57.145 63.365 57.655 63.390 ;
        RECT 62.385 47.480 62.955 47.505 ;
        RECT 59.890 46.960 62.955 47.480 ;
        RECT 62.385 46.935 62.955 46.960 ;
      LAYER met4 ;
        RECT -327.460 427.570 -322.290 427.630 ;
        RECT -321.825 427.570 -292.215 442.115 ;
        RECT -290.225 427.570 -260.615 442.115 ;
        RECT -258.625 427.570 -229.015 442.115 ;
        RECT -227.025 427.570 -197.415 442.115 ;
        RECT -195.425 427.570 -165.815 442.115 ;
        RECT -163.825 427.570 -134.215 442.115 ;
        RECT -132.225 427.570 -102.615 442.115 ;
        RECT -100.625 427.570 -71.015 442.115 ;
        RECT -69.025 427.570 -39.415 442.115 ;
        RECT -37.425 427.570 -7.815 442.115 ;
        RECT -5.825 427.570 23.785 442.115 ;
        RECT 25.775 427.570 55.385 442.115 ;
        RECT -327.460 427.110 56.380 427.570 ;
        RECT -327.460 394.510 -326.940 427.110 ;
        RECT -322.820 427.050 56.380 427.110 ;
        RECT -321.825 412.505 -292.215 427.050 ;
        RECT -290.225 412.505 -260.615 427.050 ;
        RECT -258.625 412.505 -229.015 427.050 ;
        RECT -227.025 412.505 -197.415 427.050 ;
        RECT -195.425 412.505 -165.815 427.050 ;
        RECT -163.825 412.505 -134.215 427.050 ;
        RECT -132.225 412.505 -102.615 427.050 ;
        RECT -100.625 412.505 -71.015 427.050 ;
        RECT -69.025 412.505 -39.415 427.050 ;
        RECT -37.425 412.505 -7.815 427.050 ;
        RECT -5.825 412.505 23.785 427.050 ;
        RECT 25.775 412.505 55.385 427.050 ;
        RECT -322.820 411.110 56.380 411.170 ;
        RECT -324.780 410.650 56.380 411.110 ;
        RECT -324.780 410.590 -322.380 410.650 ;
        RECT -324.780 395.725 -324.260 410.590 ;
        RECT -324.785 395.195 -324.255 395.725 ;
        RECT -321.825 394.510 -292.215 409.055 ;
        RECT -290.225 394.510 -260.615 409.055 ;
        RECT -258.625 394.510 -229.015 409.055 ;
        RECT -227.025 394.510 -197.415 409.055 ;
        RECT -195.425 394.510 -165.815 409.055 ;
        RECT -163.825 394.510 -134.215 409.055 ;
        RECT -132.225 394.510 -102.615 409.055 ;
        RECT -100.625 394.510 -71.015 409.055 ;
        RECT -69.025 394.510 -39.415 409.055 ;
        RECT -37.425 394.510 -7.815 409.055 ;
        RECT -5.825 394.510 23.785 409.055 ;
        RECT 25.775 394.510 55.385 409.055 ;
        RECT -327.460 394.490 56.380 394.510 ;
        RECT -327.460 393.990 59.910 394.490 ;
        RECT -324.780 378.110 -324.260 392.790 ;
        RECT -321.825 379.445 -292.215 393.990 ;
        RECT -290.225 379.445 -260.615 393.990 ;
        RECT -258.625 379.445 -229.015 393.990 ;
        RECT -227.025 379.445 -197.415 393.990 ;
        RECT -195.425 379.445 -165.815 393.990 ;
        RECT -163.825 379.445 -134.215 393.990 ;
        RECT -132.225 379.445 -102.615 393.990 ;
        RECT -100.625 379.445 -71.015 393.990 ;
        RECT -69.025 379.445 -39.415 393.990 ;
        RECT -37.425 379.445 -7.815 393.990 ;
        RECT -5.825 379.445 23.785 393.990 ;
        RECT 25.775 379.445 55.385 393.990 ;
        RECT 55.920 393.970 59.910 393.990 ;
        RECT -324.780 378.085 56.380 378.110 ;
        RECT -324.780 377.590 57.325 378.085 ;
        RECT 55.915 377.555 57.325 377.590 ;
        RECT -321.825 361.450 -292.215 375.995 ;
        RECT -290.225 361.450 -260.615 375.995 ;
        RECT -258.625 361.450 -229.015 375.995 ;
        RECT -227.025 361.450 -197.415 375.995 ;
        RECT -195.425 361.450 -165.815 375.995 ;
        RECT -163.825 361.450 -134.215 375.995 ;
        RECT -132.225 361.450 -102.615 375.995 ;
        RECT -100.625 361.450 -71.015 375.995 ;
        RECT -69.025 361.450 -39.415 375.995 ;
        RECT -37.425 361.450 -7.815 375.995 ;
        RECT -5.825 361.450 23.785 375.995 ;
        RECT 25.775 361.450 55.385 375.995 ;
        RECT 56.795 362.225 57.325 377.555 ;
        RECT 59.390 361.450 59.910 393.970 ;
        RECT -322.820 361.400 59.910 361.450 ;
        RECT -326.020 360.930 59.910 361.400 ;
        RECT -326.020 360.880 -322.250 360.930 ;
        RECT -326.020 328.390 -325.500 360.880 ;
        RECT -321.825 346.385 -292.215 360.930 ;
        RECT -290.225 346.385 -260.615 360.930 ;
        RECT -258.625 346.385 -229.015 360.930 ;
        RECT -227.025 346.385 -197.415 360.930 ;
        RECT -195.425 346.385 -165.815 360.930 ;
        RECT -163.825 346.385 -134.215 360.930 ;
        RECT -132.225 346.385 -102.615 360.930 ;
        RECT -100.625 346.385 -71.015 360.930 ;
        RECT -69.025 346.385 -39.415 360.930 ;
        RECT -37.425 346.385 -7.815 360.930 ;
        RECT -5.825 346.385 23.785 360.930 ;
        RECT 25.775 346.385 55.385 360.930 ;
        RECT 56.800 345.050 57.320 359.730 ;
        RECT -322.820 345.010 57.320 345.050 ;
        RECT -323.910 344.530 57.320 345.010 ;
        RECT -323.910 344.490 -322.230 344.530 ;
        RECT -323.910 329.255 -323.390 344.490 ;
        RECT -323.915 328.725 -323.385 329.255 ;
        RECT -321.825 328.390 -292.215 342.935 ;
        RECT -290.225 328.390 -260.615 342.935 ;
        RECT -258.625 328.390 -229.015 342.935 ;
        RECT -227.025 328.390 -197.415 342.935 ;
        RECT -195.425 328.390 -165.815 342.935 ;
        RECT -163.825 328.390 -134.215 342.935 ;
        RECT -132.225 328.390 -102.615 342.935 ;
        RECT -100.625 328.390 -71.015 342.935 ;
        RECT -69.025 328.390 -39.415 342.935 ;
        RECT -37.425 328.390 -7.815 342.935 ;
        RECT -5.825 328.390 23.785 342.935 ;
        RECT 25.775 328.390 55.385 342.935 ;
        RECT -326.020 328.350 56.380 328.390 ;
        RECT -326.020 327.870 61.220 328.350 ;
        RECT -323.910 311.990 -323.390 327.010 ;
        RECT -321.825 313.325 -292.215 327.870 ;
        RECT -290.225 313.325 -260.615 327.870 ;
        RECT -258.625 313.325 -229.015 327.870 ;
        RECT -227.025 313.325 -197.415 327.870 ;
        RECT -195.425 313.325 -165.815 327.870 ;
        RECT -163.825 313.325 -134.215 327.870 ;
        RECT -132.225 313.325 -102.615 327.870 ;
        RECT -100.625 313.325 -71.015 327.870 ;
        RECT -69.025 313.325 -39.415 327.870 ;
        RECT -37.425 313.325 -7.815 327.870 ;
        RECT -5.825 313.325 23.785 327.870 ;
        RECT 25.775 313.325 55.385 327.870 ;
        RECT 56.030 327.830 61.220 327.870 ;
        RECT 55.810 311.990 57.370 312.040 ;
        RECT -323.910 311.520 57.370 311.990 ;
        RECT -323.910 311.470 56.380 311.520 ;
        RECT -325.290 295.330 -322.250 295.420 ;
        RECT -321.825 295.330 -292.215 309.875 ;
        RECT -290.225 295.330 -260.615 309.875 ;
        RECT -258.625 295.330 -229.015 309.875 ;
        RECT -227.025 295.330 -197.415 309.875 ;
        RECT -195.425 295.330 -165.815 309.875 ;
        RECT -163.825 295.330 -134.215 309.875 ;
        RECT -132.225 295.330 -102.615 309.875 ;
        RECT -100.625 295.330 -71.015 309.875 ;
        RECT -69.025 295.330 -39.415 309.875 ;
        RECT -37.425 295.330 -7.815 309.875 ;
        RECT -5.825 295.330 23.785 309.875 ;
        RECT 25.775 295.330 55.385 309.875 ;
        RECT 56.850 297.235 57.370 311.520 ;
        RECT 56.845 296.705 57.375 297.235 ;
        RECT 60.700 295.330 61.220 327.830 ;
        RECT -325.290 294.900 61.220 295.330 ;
        RECT -325.290 262.270 -324.770 294.900 ;
        RECT -322.820 294.810 61.220 294.900 ;
        RECT -321.825 280.265 -292.215 294.810 ;
        RECT -290.225 280.265 -260.615 294.810 ;
        RECT -258.625 280.265 -229.015 294.810 ;
        RECT -227.025 280.265 -197.415 294.810 ;
        RECT -195.425 280.265 -165.815 294.810 ;
        RECT -163.825 280.265 -134.215 294.810 ;
        RECT -132.225 280.265 -102.615 294.810 ;
        RECT -100.625 280.265 -71.015 294.810 ;
        RECT -69.025 280.265 -39.415 294.810 ;
        RECT -37.425 280.265 -7.815 294.810 ;
        RECT -5.825 280.265 23.785 294.810 ;
        RECT 25.775 280.265 55.385 294.810 ;
        RECT 56.850 278.930 57.370 293.930 ;
        RECT -322.820 278.830 57.370 278.930 ;
        RECT -324.060 278.410 57.370 278.830 ;
        RECT -324.060 278.310 -322.410 278.410 ;
        RECT -324.060 263.275 -323.540 278.310 ;
        RECT -324.065 262.745 -323.535 263.275 ;
        RECT -321.825 262.270 -292.215 276.815 ;
        RECT -290.225 262.270 -260.615 276.815 ;
        RECT -258.625 262.270 -229.015 276.815 ;
        RECT -227.025 262.270 -197.415 276.815 ;
        RECT -195.425 262.270 -165.815 276.815 ;
        RECT -163.825 262.270 -134.215 276.815 ;
        RECT -132.225 262.270 -102.615 276.815 ;
        RECT -100.625 262.270 -71.015 276.815 ;
        RECT -69.025 262.270 -39.415 276.815 ;
        RECT -37.425 262.270 -7.815 276.815 ;
        RECT -5.825 262.270 23.785 276.815 ;
        RECT 25.775 262.270 55.385 276.815 ;
        RECT 55.870 262.270 60.480 262.310 ;
        RECT -325.290 261.790 60.480 262.270 ;
        RECT -325.290 261.750 56.380 261.790 ;
        RECT -324.060 245.870 -323.540 260.880 ;
        RECT -321.825 247.205 -292.215 261.750 ;
        RECT -290.225 247.205 -260.615 261.750 ;
        RECT -258.625 247.205 -229.015 261.750 ;
        RECT -227.025 247.205 -197.415 261.750 ;
        RECT -195.425 247.205 -165.815 261.750 ;
        RECT -163.825 247.205 -134.215 261.750 ;
        RECT -132.225 247.205 -102.615 261.750 ;
        RECT -100.625 247.205 -71.015 261.750 ;
        RECT -69.025 247.205 -39.415 261.750 ;
        RECT -37.425 247.205 -7.815 261.750 ;
        RECT -5.825 247.205 23.785 261.750 ;
        RECT 25.775 247.205 55.385 261.750 ;
        RECT 56.040 245.870 57.410 245.910 ;
        RECT -324.060 245.390 57.410 245.870 ;
        RECT -324.060 245.350 56.380 245.390 ;
        RECT -321.825 229.210 -292.215 243.755 ;
        RECT -290.225 229.210 -260.615 243.755 ;
        RECT -258.625 229.210 -229.015 243.755 ;
        RECT -227.025 229.210 -197.415 243.755 ;
        RECT -195.425 229.210 -165.815 243.755 ;
        RECT -163.825 229.210 -134.215 243.755 ;
        RECT -132.225 229.210 -102.615 243.755 ;
        RECT -100.625 229.210 -71.015 243.755 ;
        RECT -69.025 229.210 -39.415 243.755 ;
        RECT -37.425 229.210 -7.815 243.755 ;
        RECT -5.825 229.210 23.785 243.755 ;
        RECT 25.775 229.210 55.385 243.755 ;
        RECT 56.890 230.425 57.410 245.390 ;
        RECT 56.885 229.895 57.415 230.425 ;
        RECT 59.960 229.210 60.480 261.790 ;
        RECT -327.630 228.690 60.480 229.210 ;
        RECT -327.630 196.150 -327.110 228.690 ;
        RECT -321.825 214.145 -292.215 228.690 ;
        RECT -290.225 214.145 -260.615 228.690 ;
        RECT -258.625 214.145 -229.015 228.690 ;
        RECT -227.025 214.145 -197.415 228.690 ;
        RECT -195.425 214.145 -165.815 228.690 ;
        RECT -163.825 214.145 -134.215 228.690 ;
        RECT -132.225 214.145 -102.615 228.690 ;
        RECT -100.625 214.145 -71.015 228.690 ;
        RECT -69.025 214.145 -39.415 228.690 ;
        RECT -37.425 214.145 -7.815 228.690 ;
        RECT -5.825 214.145 23.785 228.690 ;
        RECT 25.775 214.145 55.385 228.690 ;
        RECT -324.460 212.810 -321.900 212.840 ;
        RECT 56.890 212.810 57.410 227.690 ;
        RECT 96.055 214.325 96.600 214.330 ;
        RECT -324.460 212.320 57.410 212.810 ;
        RECT -324.460 197.355 -323.940 212.320 ;
        RECT -322.820 212.290 57.410 212.320 ;
        RECT -324.465 196.825 -323.935 197.355 ;
        RECT -321.825 196.150 -292.215 210.695 ;
        RECT -290.225 196.150 -260.615 210.695 ;
        RECT -258.625 196.150 -229.015 210.695 ;
        RECT -227.025 196.150 -197.415 210.695 ;
        RECT -195.425 196.150 -165.815 210.695 ;
        RECT -163.825 196.150 -134.215 210.695 ;
        RECT -132.225 196.150 -102.615 210.695 ;
        RECT -100.625 196.150 -71.015 210.695 ;
        RECT -69.025 196.150 -39.415 210.695 ;
        RECT -37.425 196.150 -7.815 210.695 ;
        RECT -5.825 196.150 23.785 210.695 ;
        RECT 25.775 196.150 55.385 210.695 ;
        RECT 55.910 196.150 58.930 196.160 ;
        RECT -327.630 195.640 58.930 196.150 ;
        RECT -327.630 195.630 56.380 195.640 ;
        RECT -324.460 179.750 -323.940 194.810 ;
        RECT -321.825 181.085 -292.215 195.630 ;
        RECT -290.225 181.085 -260.615 195.630 ;
        RECT -258.625 181.085 -229.015 195.630 ;
        RECT -227.025 181.085 -197.415 195.630 ;
        RECT -195.425 181.085 -165.815 195.630 ;
        RECT -163.825 181.085 -134.215 195.630 ;
        RECT -132.225 181.085 -102.615 195.630 ;
        RECT -100.625 181.085 -71.015 195.630 ;
        RECT -69.025 181.085 -39.415 195.630 ;
        RECT -37.425 181.085 -7.815 195.630 ;
        RECT -5.825 181.085 23.785 195.630 ;
        RECT 25.775 181.085 55.385 195.630 ;
        RECT -324.460 179.690 56.380 179.750 ;
        RECT -324.460 179.230 57.600 179.690 ;
        RECT 56.170 179.170 57.600 179.230 ;
        RECT -321.825 163.090 -292.215 177.635 ;
        RECT -290.225 163.090 -260.615 177.635 ;
        RECT -258.625 163.090 -229.015 177.635 ;
        RECT -227.025 163.090 -197.415 177.635 ;
        RECT -195.425 163.090 -165.815 177.635 ;
        RECT -163.825 163.090 -134.215 177.635 ;
        RECT -132.225 163.090 -102.615 177.635 ;
        RECT -100.625 163.090 -71.015 177.635 ;
        RECT -69.025 163.090 -39.415 177.635 ;
        RECT -37.425 163.090 -7.815 177.635 ;
        RECT -5.825 163.090 23.785 177.635 ;
        RECT 25.775 163.090 55.385 177.635 ;
        RECT 57.080 164.315 57.600 179.170 ;
        RECT 57.075 163.785 57.605 164.315 ;
        RECT 58.410 163.090 58.930 195.640 ;
        RECT 92.755 181.260 93.290 214.325 ;
        RECT 96.055 214.320 97.695 214.325 ;
        RECT 96.055 213.800 255.230 214.320 ;
        RECT 96.055 213.790 97.695 213.800 ;
        RECT 96.055 213.785 96.600 213.790 ;
        RECT 254.935 181.260 258.440 181.265 ;
        RECT 92.755 180.750 258.440 181.260 ;
        RECT 92.755 180.740 255.230 180.750 ;
        RECT 92.755 180.735 93.290 180.740 ;
        RECT -322.820 163.030 58.930 163.090 ;
        RECT -326.150 162.570 58.930 163.030 ;
        RECT -326.150 162.510 -322.270 162.570 ;
        RECT -326.150 130.030 -325.630 162.510 ;
        RECT -321.825 148.025 -292.215 162.570 ;
        RECT -290.225 148.025 -260.615 162.570 ;
        RECT -258.625 148.025 -229.015 162.570 ;
        RECT -227.025 148.025 -197.415 162.570 ;
        RECT -195.425 148.025 -165.815 162.570 ;
        RECT -163.825 148.025 -134.215 162.570 ;
        RECT -132.225 148.025 -102.615 162.570 ;
        RECT -100.625 148.025 -71.015 162.570 ;
        RECT -69.025 148.025 -39.415 162.570 ;
        RECT -37.425 148.025 -7.815 162.570 ;
        RECT -5.825 148.025 23.785 162.570 ;
        RECT 25.775 148.025 55.385 162.570 ;
        RECT -324.240 146.690 -322.400 146.720 ;
        RECT 57.080 146.690 57.600 161.770 ;
        RECT 257.925 148.200 258.440 180.750 ;
        RECT 97.230 148.150 258.440 148.200 ;
        RECT -324.240 146.200 57.600 146.690 ;
        RECT -324.240 131.225 -323.720 146.200 ;
        RECT -322.820 146.170 57.600 146.200 ;
        RECT 95.640 147.680 258.440 148.150 ;
        RECT 95.640 147.630 97.560 147.680 ;
        RECT -324.245 130.695 -323.715 131.225 ;
        RECT -321.825 130.030 -292.215 144.575 ;
        RECT -290.225 130.030 -260.615 144.575 ;
        RECT -258.625 130.030 -229.015 144.575 ;
        RECT -227.025 130.030 -197.415 144.575 ;
        RECT -195.425 130.030 -165.815 144.575 ;
        RECT -163.825 130.030 -134.215 144.575 ;
        RECT -132.225 130.030 -102.615 144.575 ;
        RECT -100.625 130.030 -71.015 144.575 ;
        RECT -69.025 130.030 -39.415 144.575 ;
        RECT -37.425 130.030 -7.815 144.575 ;
        RECT -5.825 130.030 23.785 144.575 ;
        RECT 25.775 130.030 55.385 144.575 ;
        RECT 95.640 133.055 96.160 147.630 ;
        RECT 95.635 132.525 96.165 133.055 ;
        RECT -326.150 129.960 56.380 130.030 ;
        RECT -326.150 129.510 59.930 129.960 ;
        RECT -324.240 113.630 -323.720 128.740 ;
        RECT -321.825 114.965 -292.215 129.510 ;
        RECT -290.225 114.965 -260.615 129.510 ;
        RECT -258.625 114.965 -229.015 129.510 ;
        RECT -227.025 114.965 -197.415 129.510 ;
        RECT -195.425 114.965 -165.815 129.510 ;
        RECT -163.825 114.965 -134.215 129.510 ;
        RECT -132.225 114.965 -102.615 129.510 ;
        RECT -100.625 114.965 -71.015 129.510 ;
        RECT -69.025 114.965 -39.415 129.510 ;
        RECT -37.425 114.965 -7.815 129.510 ;
        RECT -5.825 114.965 23.785 129.510 ;
        RECT 25.775 114.965 55.385 129.510 ;
        RECT 56.030 129.440 59.930 129.510 ;
        RECT 55.930 113.630 57.640 113.720 ;
        RECT -324.240 113.200 57.640 113.630 ;
        RECT -324.240 113.110 56.380 113.200 ;
        RECT -321.825 96.970 -292.215 111.515 ;
        RECT -290.225 96.970 -260.615 111.515 ;
        RECT -258.625 96.970 -229.015 111.515 ;
        RECT -227.025 96.970 -197.415 111.515 ;
        RECT -195.425 96.970 -165.815 111.515 ;
        RECT -163.825 96.970 -134.215 111.515 ;
        RECT -132.225 96.970 -102.615 111.515 ;
        RECT -100.625 96.970 -71.015 111.515 ;
        RECT -69.025 96.970 -39.415 111.515 ;
        RECT -37.425 96.970 -7.815 111.515 ;
        RECT -5.825 96.970 23.785 111.515 ;
        RECT 25.775 96.970 55.385 111.515 ;
        RECT 57.120 98.025 57.640 113.200 ;
        RECT 57.115 97.495 57.645 98.025 ;
        RECT 59.410 96.970 59.930 129.440 ;
        RECT 95.640 115.140 96.160 129.980 ;
        RECT 255.625 115.160 256.155 115.165 ;
        RECT 254.680 115.140 256.155 115.160 ;
        RECT 95.640 114.640 256.155 115.140 ;
        RECT 95.640 114.620 255.230 114.640 ;
        RECT 255.625 114.635 256.155 114.640 ;
        RECT -322.820 96.820 59.930 96.970 ;
        RECT -326.940 96.450 59.930 96.820 ;
        RECT -326.940 96.300 -322.350 96.450 ;
        RECT -326.940 63.910 -326.420 96.300 ;
        RECT -321.825 81.905 -292.215 96.450 ;
        RECT -290.225 81.905 -260.615 96.450 ;
        RECT -258.625 81.905 -229.015 96.450 ;
        RECT -227.025 81.905 -197.415 96.450 ;
        RECT -195.425 81.905 -165.815 96.450 ;
        RECT -163.825 81.905 -134.215 96.450 ;
        RECT -132.225 81.905 -102.615 96.450 ;
        RECT -100.625 81.905 -71.015 96.450 ;
        RECT -69.025 81.905 -39.415 96.450 ;
        RECT -37.425 81.905 -7.815 96.450 ;
        RECT -5.825 81.905 23.785 96.450 ;
        RECT 25.775 81.905 55.385 96.450 ;
        RECT -325.110 80.570 -322.190 80.620 ;
        RECT 57.120 80.570 57.640 95.700 ;
        RECT 82.915 87.700 83.445 87.705 ;
        RECT 82.915 87.180 96.130 87.700 ;
        RECT 82.915 87.175 83.445 87.180 ;
        RECT 95.610 82.060 96.130 87.180 ;
        RECT 258.290 82.080 258.810 115.160 ;
        RECT 97.230 82.060 258.810 82.080 ;
        RECT 95.610 81.560 258.810 82.060 ;
        RECT 95.610 81.540 97.680 81.560 ;
        RECT -325.110 80.100 57.640 80.570 ;
        RECT -325.110 65.975 -324.590 80.100 ;
        RECT -322.820 80.050 57.640 80.100 ;
        RECT -325.115 65.445 -324.585 65.975 ;
        RECT -321.825 63.910 -292.215 78.455 ;
        RECT -290.225 63.910 -260.615 78.455 ;
        RECT -258.625 63.910 -229.015 78.455 ;
        RECT -227.025 63.910 -197.415 78.455 ;
        RECT -195.425 63.910 -165.815 78.455 ;
        RECT -163.825 63.910 -134.215 78.455 ;
        RECT -132.225 63.910 -102.615 78.455 ;
        RECT -100.625 63.910 -71.015 78.455 ;
        RECT -69.025 63.910 -39.415 78.455 ;
        RECT -37.425 63.910 -7.815 78.455 ;
        RECT -5.825 63.910 23.785 78.455 ;
        RECT 25.775 63.910 55.385 78.455 ;
        RECT -326.940 63.390 57.660 63.910 ;
        RECT -325.110 47.510 -324.590 62.400 ;
        RECT -321.825 48.845 -292.215 63.390 ;
        RECT -290.225 48.845 -260.615 63.390 ;
        RECT -258.625 48.845 -229.015 63.390 ;
        RECT -227.025 48.845 -197.415 63.390 ;
        RECT -195.425 48.845 -165.815 63.390 ;
        RECT -163.825 48.845 -134.215 63.390 ;
        RECT -132.225 48.845 -102.615 63.390 ;
        RECT -100.625 48.845 -71.015 63.390 ;
        RECT -69.025 48.845 -39.415 63.390 ;
        RECT -37.425 48.845 -7.815 63.390 ;
        RECT -5.825 48.845 23.785 63.390 ;
        RECT 25.775 48.845 55.385 63.390 ;
        RECT -325.110 47.480 57.400 47.510 ;
        RECT 59.915 47.480 60.445 47.485 ;
        RECT -325.110 46.990 60.445 47.480 ;
        RECT 56.830 46.960 60.445 46.990 ;
        RECT 59.915 46.955 60.445 46.960 ;
  END
END cp
MACRO pll
  CLASS BLOCK ;
  FOREIGN pll ;
  ORIGIN 324.520 18.235 ;
  SIZE 586.465 BY 449.165 ;
  OBS
      LAYER pwell ;
        RECT 59.850 31.620 61.890 32.050 ;
        RECT 59.850 24.970 60.280 31.620 ;
        RECT 61.460 24.970 61.890 31.620 ;
      LAYER nwell ;
        RECT 103.975 29.230 108.665 31.340 ;
        RECT 124.325 28.510 129.015 30.620 ;
        RECT 152.910 28.860 157.600 30.970 ;
      LAYER pwell ;
        RECT 104.855 26.440 107.855 28.450 ;
      LAYER nwell ;
        RECT 173.260 28.140 177.950 30.250 ;
      LAYER pwell ;
        RECT 125.045 25.690 128.045 27.700 ;
        RECT 153.790 26.070 156.790 28.080 ;
        RECT 173.980 25.320 176.980 27.330 ;
        RECT 59.850 24.540 61.890 24.970 ;
      LAYER nwell ;
        RECT -2.680 20.450 44.510 22.590 ;
        RECT 90.640 17.890 92.750 22.580 ;
        RECT 94.665 18.320 99.355 20.430 ;
        RECT 104.145 17.690 106.255 22.380 ;
        RECT 109.595 17.680 111.705 22.370 ;
        RECT 114.365 18.800 119.055 20.910 ;
        RECT 4.390 13.920 6.530 16.650 ;
        RECT -28.260 10.915 -7.180 12.520 ;
      LAYER pwell ;
        RECT 4.460 11.240 6.500 13.660 ;
      LAYER nwell ;
        RECT 12.520 12.510 14.660 16.700 ;
        RECT 22.830 13.720 24.970 16.450 ;
        RECT 28.540 13.840 30.680 16.570 ;
      LAYER pwell ;
        RECT 90.670 14.310 92.680 17.310 ;
        RECT 95.455 15.510 98.455 17.520 ;
        RECT 104.225 14.520 106.235 17.520 ;
        RECT 109.705 14.140 111.715 17.140 ;
        RECT 115.255 16.090 118.255 18.100 ;
      LAYER nwell ;
        RECT 122.955 18.050 125.065 22.740 ;
        RECT 127.975 17.820 130.085 22.510 ;
      LAYER pwell ;
        RECT 123.035 14.780 125.045 17.780 ;
      LAYER nwell ;
        RECT 139.575 17.520 141.685 22.210 ;
        RECT 143.600 17.950 148.290 20.060 ;
      LAYER pwell ;
        RECT 128.055 14.480 130.065 17.480 ;
      LAYER nwell ;
        RECT 153.080 17.320 155.190 22.010 ;
        RECT 158.530 17.310 160.640 22.000 ;
        RECT 163.300 18.430 167.990 20.540 ;
      LAYER pwell ;
        RECT 139.605 13.940 141.615 16.940 ;
        RECT 144.390 15.140 147.390 17.150 ;
        RECT 153.160 14.150 155.170 17.150 ;
        RECT 158.640 13.770 160.650 16.770 ;
        RECT 164.190 15.720 167.190 17.730 ;
      LAYER nwell ;
        RECT 171.890 17.680 174.000 22.370 ;
        RECT 176.910 17.450 179.020 22.140 ;
      LAYER pwell ;
        RECT 171.970 14.410 173.980 17.410 ;
        RECT 176.990 14.110 179.000 17.110 ;
      LAYER nwell ;
        RECT 12.460 12.500 14.660 12.510 ;
        RECT 10.710 11.070 16.520 12.500 ;
      LAYER pwell ;
        RECT -27.860 9.715 -26.930 10.625 ;
        RECT -24.365 9.715 -23.015 10.625 ;
        RECT -20.040 9.715 -19.110 10.625 ;
        RECT -16.820 9.715 -15.890 10.625 ;
        RECT -13.345 9.715 -11.515 10.625 ;
        RECT -9.000 9.715 -8.070 10.625 ;
        RECT -7.815 9.800 -7.385 10.585 ;
        RECT -27.860 9.695 -27.755 9.715 ;
        RECT -27.925 9.525 -27.755 9.695 ;
        RECT -24.250 9.525 -24.080 9.715 ;
        RECT -20.040 9.695 -19.935 9.715 ;
        RECT -16.820 9.695 -16.715 9.715 ;
        RECT -20.105 9.525 -19.935 9.695 ;
        RECT -16.885 9.525 -16.715 9.695 ;
        RECT -13.200 9.525 -13.030 9.715 ;
        RECT -9.000 9.695 -8.895 9.715 ;
        RECT -9.065 9.525 -8.895 9.695 ;
        RECT -25.100 8.555 -24.930 8.745 ;
        RECT -21.250 8.605 -21.080 8.795 ;
        RECT -25.865 7.665 -25.435 8.450 ;
        RECT -25.215 7.645 -23.865 8.555 ;
        RECT -21.365 7.695 -20.015 8.605 ;
      LAYER nwell ;
        RECT 10.710 8.500 12.140 11.070 ;
      LAYER pwell ;
        RECT 12.590 8.580 14.630 11.000 ;
      LAYER nwell ;
        RECT 15.090 8.500 16.520 11.070 ;
        RECT -21.580 7.355 -19.820 7.405 ;
        RECT -25.430 7.350 -23.400 7.355 ;
        RECT -22.130 7.350 -19.820 7.355 ;
        RECT -25.430 7.335 -19.820 7.350 ;
        RECT -26.070 5.800 -19.820 7.335 ;
        RECT 10.710 7.070 16.520 8.500 ;
        RECT -26.070 5.750 -21.120 5.800 ;
        RECT -26.070 5.730 -25.230 5.750 ;
        RECT -14.800 5.105 -11.040 6.710 ;
        RECT 20.650 6.350 22.790 9.080 ;
      LAYER pwell ;
        RECT -14.605 3.905 -12.315 4.815 ;
        RECT -11.675 3.990 -11.245 4.775 ;
        RECT -14.460 3.715 -14.290 3.905 ;
      LAYER nwell ;
        RECT 5.050 0.120 7.190 2.850 ;
        RECT -6.810 -0.400 -5.970 -0.390 ;
        RECT -27.340 -1.995 -5.970 -0.400 ;
        RECT -27.340 -2.005 -6.720 -1.995 ;
      LAYER pwell ;
        RECT -26.940 -3.205 -26.010 -2.295 ;
        RECT -23.445 -3.205 -22.095 -2.295 ;
        RECT -19.120 -3.205 -18.190 -2.295 ;
        RECT -15.900 -3.205 -14.970 -2.295 ;
        RECT -12.425 -3.205 -10.595 -2.295 ;
        RECT -8.080 -3.205 -7.150 -2.295 ;
        RECT -6.605 -3.110 -6.175 -2.325 ;
        RECT 4.990 -3.100 7.030 -0.680 ;
      LAYER nwell ;
        RECT 13.410 -2.080 15.550 2.920 ;
      LAYER pwell ;
        RECT 25.930 0.900 27.970 3.320 ;
      LAYER nwell ;
        RECT 34.420 2.600 40.230 4.030 ;
      LAYER pwell ;
        RECT 119.815 3.825 121.825 6.825 ;
        RECT 124.835 3.525 126.845 6.525 ;
      LAYER nwell ;
        RECT 34.420 0.030 35.850 2.600 ;
      LAYER pwell ;
        RECT 36.330 0.120 38.370 2.540 ;
      LAYER nwell ;
        RECT 38.800 0.030 40.230 2.600 ;
      LAYER pwell ;
        RECT -26.940 -3.225 -26.835 -3.205 ;
        RECT -27.005 -3.395 -26.835 -3.225 ;
        RECT -23.330 -3.395 -23.160 -3.205 ;
        RECT -19.120 -3.225 -19.015 -3.205 ;
        RECT -15.900 -3.225 -15.795 -3.205 ;
        RECT -19.185 -3.395 -19.015 -3.225 ;
        RECT -15.965 -3.395 -15.795 -3.225 ;
        RECT -12.280 -3.395 -12.110 -3.205 ;
        RECT -8.080 -3.225 -7.975 -3.205 ;
        RECT -8.145 -3.395 -7.975 -3.225 ;
      LAYER nwell ;
        RECT 11.770 -3.510 17.580 -2.080 ;
      LAYER pwell ;
        RECT -22.860 -3.805 -22.690 -3.615 ;
        RECT -23.925 -4.715 -22.575 -3.805 ;
        RECT -19.630 -3.865 -19.460 -3.675 ;
        RECT -20.695 -4.775 -19.345 -3.865 ;
        RECT -19.095 -4.805 -18.665 -4.020 ;
      LAYER nwell ;
        RECT -24.120 -5.065 -20.150 -5.005 ;
        RECT -24.120 -5.135 -19.130 -5.065 ;
        RECT -24.120 -6.610 -18.460 -5.135 ;
        RECT -20.890 -6.670 -18.460 -6.610 ;
        RECT -19.300 -6.740 -18.460 -6.670 ;
        RECT 11.770 -6.080 13.200 -3.510 ;
      LAYER pwell ;
        RECT 13.570 -6.020 15.610 -3.600 ;
      LAYER nwell ;
        RECT 16.150 -6.080 17.580 -3.510 ;
        RECT 11.770 -7.510 17.580 -6.080 ;
        RECT 23.090 -2.200 28.900 -0.770 ;
        RECT 34.420 -1.400 40.230 0.030 ;
        RECT 23.090 -4.770 24.520 -2.200 ;
      LAYER pwell ;
        RECT 25.030 -4.710 27.070 -2.290 ;
      LAYER nwell ;
        RECT 27.470 -4.770 28.900 -2.200 ;
        RECT 23.090 -6.200 28.900 -4.770 ;
        RECT 48.350 -6.395 50.490 -2.405 ;
        RECT 57.110 -6.385 59.250 -0.655 ;
        RECT 64.700 -6.335 66.840 -0.605 ;
        RECT 72.310 -6.315 74.450 -0.585 ;
        RECT 80.310 -6.355 82.450 -0.625 ;
        RECT 88.120 -6.335 90.260 -0.605 ;
        RECT 95.710 -6.355 97.850 -0.625 ;
        RECT 103.100 -6.385 105.240 -0.655 ;
        RECT 119.795 -1.205 121.905 3.485 ;
        RECT 124.815 -1.435 126.925 3.255 ;
      LAYER pwell ;
        RECT 131.625 3.205 134.625 5.215 ;
        RECT 138.165 4.165 140.175 7.165 ;
        RECT 143.645 3.785 145.655 6.785 ;
        RECT 151.425 3.785 154.425 5.795 ;
        RECT 157.200 3.995 159.210 6.995 ;
      LAYER nwell ;
        RECT 130.825 0.395 135.515 2.505 ;
        RECT 138.175 -1.065 140.285 3.625 ;
        RECT 143.625 -1.075 145.735 3.615 ;
        RECT 150.525 0.875 155.215 2.985 ;
        RECT 157.130 -1.275 159.240 3.415 ;
        RECT 109.620 -5.695 111.760 -2.785 ;
      LAYER pwell ;
        RECT 48.390 -9.735 50.430 -7.315 ;
        RECT 57.170 -9.095 59.210 -6.675 ;
        RECT 64.760 -9.045 66.800 -6.625 ;
        RECT 72.370 -9.025 74.410 -6.605 ;
        RECT 17.060 -12.540 34.060 -10.500 ;
        RECT 57.180 -11.525 59.220 -9.105 ;
        RECT 64.770 -11.475 66.810 -9.055 ;
        RECT 72.380 -11.455 74.420 -9.035 ;
        RECT 80.370 -9.065 82.410 -6.645 ;
        RECT 88.180 -9.045 90.220 -6.625 ;
        RECT 80.380 -11.495 82.420 -9.075 ;
        RECT 88.190 -11.475 90.230 -9.055 ;
        RECT 95.770 -9.065 97.810 -6.645 ;
        RECT 95.780 -11.495 97.820 -9.075 ;
        RECT 103.160 -9.095 105.200 -6.675 ;
        RECT 109.620 -8.645 111.660 -6.225 ;
        RECT 121.835 -6.395 124.835 -4.385 ;
        RECT 142.025 -7.145 145.025 -5.135 ;
        RECT 103.170 -11.525 105.210 -9.105 ;
      LAYER nwell ;
        RECT 120.865 -9.315 125.555 -7.205 ;
        RECT 141.215 -10.035 145.905 -7.925 ;
      LAYER li1 ;
        RECT 59.980 31.750 61.760 31.920 ;
        RECT 59.980 24.840 60.150 31.750 ;
        RECT 60.630 31.020 61.110 31.190 ;
        RECT 60.710 29.205 61.030 31.020 ;
        RECT 60.710 25.570 61.030 27.385 ;
        RECT 60.630 25.400 61.110 25.570 ;
        RECT 61.590 24.840 61.760 31.750 ;
        RECT 104.155 30.990 108.485 31.160 ;
        RECT 104.155 29.580 104.325 30.990 ;
        RECT 108.315 30.670 108.485 30.990 ;
        RECT 104.665 30.120 104.835 30.450 ;
        RECT 105.050 30.420 107.590 30.590 ;
        RECT 105.050 29.980 107.590 30.150 ;
        RECT 107.805 30.120 107.975 30.450 ;
        RECT 108.315 29.920 108.625 30.670 ;
        RECT 153.090 30.620 157.420 30.790 ;
        RECT 124.505 30.270 128.835 30.440 ;
        RECT 108.315 29.580 108.485 29.920 ;
        RECT 104.155 29.410 108.485 29.580 ;
        RECT 124.505 28.860 124.675 30.270 ;
        RECT 125.015 29.400 125.185 29.730 ;
        RECT 125.400 29.700 127.940 29.870 ;
        RECT 125.400 29.260 127.940 29.430 ;
        RECT 128.155 29.400 128.325 29.730 ;
        RECT 128.665 28.860 128.835 30.270 ;
        RECT 153.090 29.210 153.260 30.620 ;
        RECT 157.250 30.300 157.420 30.620 ;
        RECT 153.600 29.750 153.770 30.080 ;
        RECT 153.985 30.050 156.525 30.220 ;
        RECT 153.985 29.610 156.525 29.780 ;
        RECT 156.740 29.750 156.910 30.080 ;
        RECT 157.250 29.550 157.560 30.300 ;
        RECT 173.440 29.900 177.770 30.070 ;
        RECT 157.250 29.210 157.420 29.550 ;
        RECT 153.090 29.040 157.420 29.210 ;
        RECT 124.505 28.690 128.835 28.860 ;
        RECT 173.440 28.490 173.610 29.900 ;
        RECT 173.950 29.030 174.120 29.360 ;
        RECT 174.335 29.330 176.875 29.500 ;
        RECT 174.335 28.890 176.875 29.060 ;
        RECT 177.090 29.030 177.260 29.360 ;
        RECT 177.600 28.490 177.770 29.900 ;
        RECT 173.440 28.320 177.770 28.490 ;
        RECT 104.985 28.150 107.725 28.320 ;
        RECT 104.985 27.910 105.155 28.150 ;
        RECT 104.785 27.010 105.155 27.910 ;
        RECT 105.495 27.280 105.665 27.610 ;
        RECT 105.835 27.580 106.875 27.750 ;
        RECT 105.835 27.140 106.875 27.310 ;
        RECT 107.045 27.280 107.215 27.610 ;
        RECT 104.985 26.740 105.155 27.010 ;
        RECT 107.555 26.740 107.725 28.150 ;
        RECT 153.920 27.780 156.660 27.950 ;
        RECT 125.175 27.400 127.915 27.570 ;
        RECT 153.920 27.540 154.090 27.780 ;
        RECT 125.175 27.180 125.345 27.400 ;
        RECT 104.985 26.570 107.725 26.740 ;
        RECT 125.165 26.300 125.365 27.180 ;
        RECT 125.685 26.530 125.855 26.860 ;
        RECT 126.025 26.830 127.065 27.000 ;
        RECT 126.025 26.390 127.065 26.560 ;
        RECT 127.235 26.530 127.405 26.860 ;
        RECT 125.175 25.990 125.345 26.300 ;
        RECT 127.745 25.990 127.915 27.400 ;
        RECT 153.720 26.640 154.090 27.540 ;
        RECT 154.430 26.910 154.600 27.240 ;
        RECT 154.770 27.210 155.810 27.380 ;
        RECT 154.770 26.770 155.810 26.940 ;
        RECT 155.980 26.910 156.150 27.240 ;
        RECT 153.920 26.370 154.090 26.640 ;
        RECT 156.490 26.370 156.660 27.780 ;
        RECT 174.110 27.030 176.850 27.200 ;
        RECT 174.110 26.810 174.280 27.030 ;
        RECT 153.920 26.200 156.660 26.370 ;
        RECT 125.175 25.820 127.915 25.990 ;
        RECT 174.100 25.930 174.300 26.810 ;
        RECT 174.620 26.160 174.790 26.490 ;
        RECT 174.960 26.460 176.000 26.630 ;
        RECT 174.960 26.020 176.000 26.190 ;
        RECT 176.170 26.160 176.340 26.490 ;
        RECT 174.110 25.620 174.280 25.930 ;
        RECT 176.680 25.620 176.850 27.030 ;
        RECT 174.110 25.450 176.850 25.620 ;
        RECT 59.980 24.670 61.760 24.840 ;
        RECT 123.555 22.560 124.465 22.720 ;
        RECT -2.500 22.240 44.330 22.410 ;
        RECT 91.230 22.400 92.200 22.530 ;
        RECT -2.500 20.800 -2.330 22.240 ;
        RECT -1.990 21.355 -1.820 21.685 ;
        RECT -1.605 21.670 43.435 21.840 ;
        RECT -1.605 21.200 43.435 21.370 ;
        RECT 43.650 21.355 43.820 21.685 ;
        RECT 44.160 20.800 44.330 22.240 ;
        RECT -2.500 20.630 44.330 20.800 ;
        RECT 90.820 22.230 92.570 22.400 ;
        RECT 123.135 22.390 124.885 22.560 ;
        RECT 90.820 18.240 90.990 22.230 ;
        RECT 91.530 21.720 91.860 21.890 ;
        RECT 91.390 18.965 91.560 21.505 ;
        RECT 91.830 18.965 92.000 21.505 ;
        RECT 91.530 18.580 91.860 18.750 ;
        RECT 92.400 18.240 92.570 22.230 ;
        RECT 104.745 22.200 105.685 22.240 ;
        RECT 104.325 22.030 106.075 22.200 ;
        RECT 110.105 22.190 111.075 22.330 ;
        RECT 94.845 20.080 99.175 20.250 ;
        RECT 94.845 18.670 95.015 20.080 ;
        RECT 99.005 19.820 99.175 20.080 ;
        RECT 95.355 19.210 95.525 19.540 ;
        RECT 95.740 19.510 98.280 19.680 ;
        RECT 95.740 19.070 98.280 19.240 ;
        RECT 98.495 19.210 98.665 19.540 ;
        RECT 99.005 18.970 99.240 19.820 ;
        RECT 99.005 18.670 99.175 18.970 ;
        RECT 94.845 18.500 99.175 18.670 ;
        RECT 90.820 18.070 92.570 18.240 ;
        RECT 104.325 18.040 104.495 22.030 ;
        RECT 105.035 21.520 105.365 21.690 ;
        RECT 104.895 18.765 105.065 21.305 ;
        RECT 105.335 18.765 105.505 21.305 ;
        RECT 105.035 18.380 105.365 18.550 ;
        RECT 105.905 18.040 106.075 22.030 ;
        RECT 104.325 17.870 106.075 18.040 ;
        RECT 109.775 22.020 111.525 22.190 ;
        RECT 109.775 18.030 109.945 22.020 ;
        RECT 110.485 21.510 110.815 21.680 ;
        RECT 110.345 18.755 110.515 21.295 ;
        RECT 110.785 18.755 110.955 21.295 ;
        RECT 110.485 18.370 110.815 18.540 ;
        RECT 111.355 18.030 111.525 22.020 ;
        RECT 114.545 20.560 118.875 20.730 ;
        RECT 114.545 19.150 114.715 20.560 ;
        RECT 118.705 20.420 118.875 20.560 ;
        RECT 115.055 19.690 115.225 20.020 ;
        RECT 115.440 19.990 117.980 20.160 ;
        RECT 115.440 19.550 117.980 19.720 ;
        RECT 118.195 19.690 118.365 20.020 ;
        RECT 118.705 19.310 118.985 20.420 ;
        RECT 118.705 19.150 118.875 19.310 ;
        RECT 114.545 18.980 118.875 19.150 ;
        RECT 123.135 18.400 123.305 22.390 ;
        RECT 123.555 22.380 124.465 22.390 ;
        RECT 123.845 21.880 124.175 22.050 ;
        RECT 123.705 19.125 123.875 21.665 ;
        RECT 124.145 19.125 124.315 21.665 ;
        RECT 123.845 18.740 124.175 18.910 ;
        RECT 124.715 18.400 124.885 22.390 ;
        RECT 128.560 22.330 129.530 22.480 ;
        RECT 123.135 18.230 124.885 18.400 ;
        RECT 128.155 22.160 129.905 22.330 ;
        RECT 172.490 22.190 173.400 22.350 ;
        RECT 109.775 17.860 111.525 18.030 ;
        RECT 128.155 18.170 128.325 22.160 ;
        RECT 128.865 21.650 129.195 21.820 ;
        RECT 128.725 18.895 128.895 21.435 ;
        RECT 129.165 18.895 129.335 21.435 ;
        RECT 128.865 18.510 129.195 18.680 ;
        RECT 129.735 18.170 129.905 22.160 ;
        RECT 140.165 22.030 141.135 22.160 ;
        RECT 128.155 18.000 129.905 18.170 ;
        RECT 139.755 21.860 141.505 22.030 ;
        RECT 172.070 22.020 173.820 22.190 ;
        RECT 115.385 17.800 118.125 17.970 ;
        RECT 115.385 17.640 115.555 17.800 ;
        RECT 95.585 17.220 98.325 17.390 ;
        RECT 90.800 17.010 92.550 17.180 ;
        RECT 4.570 16.300 6.350 16.470 ;
        RECT 4.570 14.270 4.740 16.300 ;
        RECT 5.295 15.790 5.625 15.960 ;
        RECT 5.140 14.995 5.310 15.575 ;
        RECT 5.610 14.995 5.780 15.575 ;
        RECT 5.295 14.610 5.625 14.780 ;
        RECT 6.180 14.270 6.350 16.300 ;
        RECT 4.570 14.100 6.350 14.270 ;
        RECT 12.700 16.350 14.480 16.520 ;
        RECT 12.700 14.320 12.870 16.350 ;
        RECT 13.425 15.840 13.755 16.010 ;
        RECT 13.270 15.045 13.440 15.625 ;
        RECT 13.740 15.045 13.910 15.625 ;
        RECT 13.425 14.660 13.755 14.830 ;
        RECT 14.310 14.320 14.480 16.350 ;
        RECT 12.700 14.150 14.480 14.320 ;
        RECT 23.010 16.100 24.790 16.270 ;
        RECT 23.010 14.070 23.180 16.100 ;
        RECT 23.735 15.590 24.065 15.760 ;
        RECT 23.580 14.795 23.750 15.375 ;
        RECT 24.050 14.795 24.220 15.375 ;
        RECT 23.735 14.410 24.065 14.580 ;
        RECT 24.620 14.070 24.790 16.100 ;
        RECT 23.010 13.900 24.790 14.070 ;
        RECT 28.720 16.220 30.500 16.390 ;
        RECT 28.720 14.190 28.890 16.220 ;
        RECT 29.445 15.710 29.775 15.880 ;
        RECT 29.290 14.915 29.460 15.495 ;
        RECT 29.760 14.915 29.930 15.495 ;
        RECT 29.445 14.530 29.775 14.700 ;
        RECT 30.330 14.190 30.500 16.220 ;
        RECT 90.800 14.610 90.970 17.010 ;
        RECT 91.510 16.500 91.840 16.670 ;
        RECT 91.370 15.290 91.540 16.330 ;
        RECT 91.810 15.290 91.980 16.330 ;
        RECT 91.510 14.950 91.840 15.120 ;
        RECT 92.380 14.610 92.550 17.010 ;
        RECT 95.585 16.980 95.755 17.220 ;
        RECT 95.500 16.120 95.755 16.980 ;
        RECT 96.095 16.350 96.265 16.680 ;
        RECT 96.435 16.650 97.475 16.820 ;
        RECT 96.435 16.210 97.475 16.380 ;
        RECT 97.645 16.350 97.815 16.680 ;
        RECT 95.585 15.810 95.755 16.120 ;
        RECT 98.155 15.810 98.325 17.220 ;
        RECT 95.585 15.640 98.325 15.810 ;
        RECT 104.355 17.220 106.105 17.390 ;
        RECT 104.355 14.820 104.525 17.220 ;
        RECT 105.065 16.710 105.395 16.880 ;
        RECT 104.925 15.500 105.095 16.540 ;
        RECT 105.365 15.500 105.535 16.540 ;
        RECT 105.065 15.160 105.395 15.330 ;
        RECT 105.935 14.820 106.105 17.220 ;
        RECT 104.355 14.650 106.105 14.820 ;
        RECT 109.835 16.840 111.585 17.010 ;
        RECT 90.800 14.440 92.550 14.610 ;
        RECT 104.795 14.580 105.665 14.650 ;
        RECT 109.835 14.440 110.005 16.840 ;
        RECT 110.545 16.330 110.875 16.500 ;
        RECT 110.405 15.120 110.575 16.160 ;
        RECT 110.845 15.120 111.015 16.160 ;
        RECT 110.545 14.780 110.875 14.950 ;
        RECT 111.415 14.440 111.585 16.840 ;
        RECT 115.325 16.670 115.555 17.640 ;
        RECT 115.895 16.930 116.065 17.260 ;
        RECT 116.235 17.230 117.275 17.400 ;
        RECT 116.235 16.790 117.275 16.960 ;
        RECT 117.445 16.930 117.615 17.260 ;
        RECT 115.385 16.390 115.555 16.670 ;
        RECT 117.955 16.390 118.125 17.800 ;
        RECT 139.755 17.870 139.925 21.860 ;
        RECT 140.465 21.350 140.795 21.520 ;
        RECT 140.325 18.595 140.495 21.135 ;
        RECT 140.765 18.595 140.935 21.135 ;
        RECT 140.465 18.210 140.795 18.380 ;
        RECT 141.335 17.870 141.505 21.860 ;
        RECT 153.680 21.830 154.620 21.870 ;
        RECT 153.260 21.660 155.010 21.830 ;
        RECT 159.040 21.820 160.010 21.960 ;
        RECT 143.780 19.710 148.110 19.880 ;
        RECT 143.780 18.300 143.950 19.710 ;
        RECT 147.940 19.450 148.110 19.710 ;
        RECT 144.290 18.840 144.460 19.170 ;
        RECT 144.675 19.140 147.215 19.310 ;
        RECT 144.675 18.700 147.215 18.870 ;
        RECT 147.430 18.840 147.600 19.170 ;
        RECT 147.940 18.600 148.175 19.450 ;
        RECT 147.940 18.300 148.110 18.600 ;
        RECT 143.780 18.130 148.110 18.300 ;
        RECT 139.755 17.700 141.505 17.870 ;
        RECT 153.260 17.670 153.430 21.660 ;
        RECT 153.970 21.150 154.300 21.320 ;
        RECT 153.830 18.395 154.000 20.935 ;
        RECT 154.270 18.395 154.440 20.935 ;
        RECT 153.970 18.010 154.300 18.180 ;
        RECT 154.840 17.670 155.010 21.660 ;
        RECT 115.385 16.220 118.125 16.390 ;
        RECT 123.165 17.480 124.915 17.650 ;
        RECT 153.260 17.500 155.010 17.670 ;
        RECT 158.710 21.650 160.460 21.820 ;
        RECT 158.710 17.660 158.880 21.650 ;
        RECT 159.420 21.140 159.750 21.310 ;
        RECT 159.280 18.385 159.450 20.925 ;
        RECT 159.720 18.385 159.890 20.925 ;
        RECT 159.420 18.000 159.750 18.170 ;
        RECT 160.290 17.660 160.460 21.650 ;
        RECT 163.480 20.190 167.810 20.360 ;
        RECT 163.480 18.780 163.650 20.190 ;
        RECT 167.640 20.050 167.810 20.190 ;
        RECT 163.990 19.320 164.160 19.650 ;
        RECT 164.375 19.620 166.915 19.790 ;
        RECT 164.375 19.180 166.915 19.350 ;
        RECT 167.130 19.320 167.300 19.650 ;
        RECT 167.640 18.940 167.920 20.050 ;
        RECT 167.640 18.780 167.810 18.940 ;
        RECT 163.480 18.610 167.810 18.780 ;
        RECT 172.070 18.030 172.240 22.020 ;
        RECT 172.490 22.010 173.400 22.020 ;
        RECT 172.780 21.510 173.110 21.680 ;
        RECT 172.640 18.755 172.810 21.295 ;
        RECT 173.080 18.755 173.250 21.295 ;
        RECT 172.780 18.370 173.110 18.540 ;
        RECT 173.650 18.030 173.820 22.020 ;
        RECT 177.495 21.960 178.465 22.110 ;
        RECT 172.070 17.860 173.820 18.030 ;
        RECT 177.090 21.790 178.840 21.960 ;
        RECT 158.710 17.490 160.460 17.660 ;
        RECT 177.090 17.800 177.260 21.790 ;
        RECT 177.800 21.280 178.130 21.450 ;
        RECT 177.660 18.525 177.830 21.065 ;
        RECT 178.100 18.525 178.270 21.065 ;
        RECT 177.800 18.140 178.130 18.310 ;
        RECT 178.670 17.800 178.840 21.790 ;
        RECT 177.090 17.630 178.840 17.800 ;
        RECT 123.165 15.080 123.335 17.480 ;
        RECT 123.875 16.970 124.205 17.140 ;
        RECT 123.735 15.760 123.905 16.800 ;
        RECT 124.175 15.760 124.345 16.800 ;
        RECT 123.875 15.420 124.205 15.590 ;
        RECT 124.745 15.080 124.915 17.480 ;
        RECT 164.320 17.430 167.060 17.600 ;
        RECT 123.165 14.910 124.915 15.080 ;
        RECT 128.185 17.180 129.935 17.350 ;
        RECT 164.320 17.270 164.490 17.430 ;
        RECT 123.620 14.830 124.450 14.910 ;
        RECT 128.185 14.780 128.355 17.180 ;
        RECT 128.895 16.670 129.225 16.840 ;
        RECT 128.755 15.460 128.925 16.500 ;
        RECT 129.195 15.460 129.365 16.500 ;
        RECT 128.895 15.120 129.225 15.290 ;
        RECT 129.765 14.780 129.935 17.180 ;
        RECT 144.520 16.850 147.260 17.020 ;
        RECT 128.185 14.610 129.935 14.780 ;
        RECT 139.735 16.640 141.485 16.810 ;
        RECT 128.620 14.490 129.480 14.610 ;
        RECT 91.250 14.380 92.100 14.440 ;
        RECT 109.835 14.270 111.585 14.440 ;
        RECT 28.720 14.020 30.500 14.190 ;
        RECT 110.160 14.160 111.250 14.270 ;
        RECT 139.735 14.240 139.905 16.640 ;
        RECT 140.445 16.130 140.775 16.300 ;
        RECT 140.305 14.920 140.475 15.960 ;
        RECT 140.745 14.920 140.915 15.960 ;
        RECT 140.445 14.580 140.775 14.750 ;
        RECT 141.315 14.240 141.485 16.640 ;
        RECT 144.520 16.610 144.690 16.850 ;
        RECT 144.435 15.750 144.690 16.610 ;
        RECT 145.030 15.980 145.200 16.310 ;
        RECT 145.370 16.280 146.410 16.450 ;
        RECT 145.370 15.840 146.410 16.010 ;
        RECT 146.580 15.980 146.750 16.310 ;
        RECT 144.520 15.440 144.690 15.750 ;
        RECT 147.090 15.440 147.260 16.850 ;
        RECT 144.520 15.270 147.260 15.440 ;
        RECT 153.290 16.850 155.040 17.020 ;
        RECT 153.290 14.450 153.460 16.850 ;
        RECT 154.000 16.340 154.330 16.510 ;
        RECT 153.860 15.130 154.030 16.170 ;
        RECT 154.300 15.130 154.470 16.170 ;
        RECT 154.000 14.790 154.330 14.960 ;
        RECT 154.870 14.450 155.040 16.850 ;
        RECT 153.290 14.280 155.040 14.450 ;
        RECT 158.770 16.470 160.520 16.640 ;
        RECT 139.735 14.070 141.485 14.240 ;
        RECT 153.730 14.210 154.600 14.280 ;
        RECT 158.770 14.070 158.940 16.470 ;
        RECT 159.480 15.960 159.810 16.130 ;
        RECT 159.340 14.750 159.510 15.790 ;
        RECT 159.780 14.750 159.950 15.790 ;
        RECT 159.480 14.410 159.810 14.580 ;
        RECT 160.350 14.070 160.520 16.470 ;
        RECT 164.260 16.300 164.490 17.270 ;
        RECT 164.830 16.560 165.000 16.890 ;
        RECT 165.170 16.860 166.210 17.030 ;
        RECT 165.170 16.420 166.210 16.590 ;
        RECT 166.380 16.560 166.550 16.890 ;
        RECT 164.320 16.020 164.490 16.300 ;
        RECT 166.890 16.020 167.060 17.430 ;
        RECT 164.320 15.850 167.060 16.020 ;
        RECT 172.100 17.110 173.850 17.280 ;
        RECT 172.100 14.710 172.270 17.110 ;
        RECT 172.810 16.600 173.140 16.770 ;
        RECT 172.670 15.390 172.840 16.430 ;
        RECT 173.110 15.390 173.280 16.430 ;
        RECT 172.810 15.050 173.140 15.220 ;
        RECT 173.680 14.710 173.850 17.110 ;
        RECT 172.100 14.540 173.850 14.710 ;
        RECT 177.120 16.810 178.870 16.980 ;
        RECT 172.555 14.460 173.385 14.540 ;
        RECT 177.120 14.410 177.290 16.810 ;
        RECT 177.830 16.300 178.160 16.470 ;
        RECT 177.690 15.090 177.860 16.130 ;
        RECT 178.130 15.090 178.300 16.130 ;
        RECT 177.830 14.750 178.160 14.920 ;
        RECT 178.700 14.410 178.870 16.810 ;
        RECT 177.120 14.240 178.870 14.410 ;
        RECT 177.555 14.120 178.415 14.240 ;
        RECT 140.185 14.010 141.035 14.070 ;
        RECT 158.770 13.900 160.520 14.070 ;
        RECT 159.095 13.790 160.185 13.900 ;
        RECT 4.590 13.360 6.370 13.530 ;
        RECT -28.070 12.245 -26.690 12.415 ;
        RECT -24.390 12.245 -23.010 12.415 ;
        RECT -20.250 12.245 -18.870 12.415 ;
        RECT -17.030 12.245 -15.650 12.415 ;
        RECT -13.350 12.245 -11.510 12.415 ;
        RECT -9.210 12.245 -7.370 12.415 ;
        RECT -27.730 11.105 -27.520 12.245 ;
        RECT -27.350 11.095 -27.020 12.075 ;
        RECT -24.305 11.105 -24.025 12.245 ;
        RECT -23.855 11.095 -23.525 12.075 ;
        RECT -23.355 11.105 -23.095 12.245 ;
        RECT -21.525 11.485 -20.775 11.740 ;
        RECT -27.750 10.910 -27.420 10.925 ;
        RECT -28.750 10.710 -27.420 10.910 ;
        RECT -27.750 10.685 -27.420 10.710 ;
        RECT -27.250 10.910 -27.020 11.095 ;
        RECT -24.295 10.910 -23.960 10.935 ;
        RECT -27.250 10.710 -23.960 10.910 ;
        RECT -27.750 9.695 -27.520 10.515 ;
        RECT -27.250 10.495 -27.020 10.710 ;
        RECT -24.295 10.665 -23.960 10.710 ;
        RECT -23.790 10.495 -23.620 11.095 ;
        RECT -23.450 10.910 -23.115 10.935 ;
        RECT -21.000 10.910 -20.810 11.485 ;
        RECT -19.910 11.105 -19.700 12.245 ;
        RECT -19.530 11.095 -19.200 12.075 ;
        RECT -16.690 11.105 -16.480 12.245 ;
        RECT -16.310 11.095 -15.980 12.075 ;
        RECT -19.930 10.910 -19.600 10.925 ;
        RECT -23.450 10.710 -22.350 10.910 ;
        RECT -21.000 10.710 -19.600 10.910 ;
        RECT -23.450 10.685 -23.115 10.710 ;
        RECT -27.350 9.865 -27.020 10.495 ;
        RECT -24.305 9.695 -23.995 10.495 ;
        RECT -23.790 10.210 -23.095 10.495 ;
        RECT -21.000 10.210 -20.800 10.710 ;
        RECT -19.930 10.685 -19.600 10.710 ;
        RECT -19.430 10.910 -19.200 11.095 ;
        RECT -16.710 10.910 -16.380 10.925 ;
        RECT -19.430 10.710 -16.380 10.910 ;
        RECT -23.790 10.010 -20.800 10.210 ;
        RECT -23.790 9.865 -23.095 10.010 ;
        RECT -19.930 9.695 -19.700 10.515 ;
        RECT -19.430 10.495 -19.200 10.710 ;
        RECT -16.710 10.685 -16.380 10.710 ;
        RECT -16.210 10.860 -15.980 11.095 ;
        RECT -14.800 10.860 -14.600 11.810 ;
        RECT -13.260 11.105 -13.005 12.245 ;
        RECT -12.835 11.275 -12.505 12.075 ;
        RECT -12.335 11.445 -12.105 12.245 ;
        RECT -11.935 11.275 -11.605 12.075 ;
        RECT -12.835 11.105 -11.605 11.275 ;
        RECT -10.300 11.260 -9.650 11.460 ;
        RECT -13.240 10.860 -13.020 10.935 ;
        RECT -16.210 10.660 -14.600 10.860 ;
        RECT -13.950 10.660 -13.020 10.860 ;
        RECT -19.530 9.865 -19.200 10.495 ;
        RECT -16.710 9.695 -16.480 10.515 ;
        RECT -16.210 10.495 -15.980 10.660 ;
        RECT -16.310 9.865 -15.980 10.495 ;
        RECT -13.950 9.810 -13.750 10.660 ;
        RECT -13.240 10.355 -13.020 10.660 ;
        RECT -12.835 10.205 -12.655 11.105 ;
        RECT -12.485 10.375 -12.110 10.935 ;
        RECT -11.905 10.910 -11.595 10.935 ;
        RECT -9.850 10.910 -9.650 11.260 ;
        RECT -8.870 11.105 -8.660 12.245 ;
        RECT -8.490 11.095 -8.160 12.075 ;
        RECT -8.890 10.910 -8.560 10.925 ;
        RECT -11.905 10.660 -10.600 10.910 ;
        RECT -9.850 10.710 -8.560 10.910 ;
        RECT -11.905 10.605 -11.595 10.660 ;
        RECT -11.935 10.205 -11.605 10.435 ;
        RECT -10.845 10.415 -10.650 10.660 ;
        RECT -13.260 9.695 -13.005 10.185 ;
        RECT -12.835 10.160 -11.605 10.205 ;
        RECT -9.850 10.160 -9.650 10.710 ;
        RECT -8.890 10.685 -8.560 10.710 ;
        RECT -8.390 10.910 -8.160 11.095 ;
        RECT -7.745 11.080 -7.455 12.245 ;
        RECT 4.590 11.540 4.760 13.360 ;
        RECT 5.315 12.850 5.645 13.020 ;
        RECT 5.160 12.220 5.330 12.680 ;
        RECT 5.630 12.220 5.800 12.680 ;
        RECT 5.315 11.880 5.645 12.050 ;
        RECT 6.200 11.540 6.370 13.360 ;
        RECT 4.590 11.370 6.370 11.540 ;
        RECT 10.995 12.045 16.235 12.215 ;
        RECT -8.390 10.710 -6.750 10.910 ;
        RECT -12.835 9.960 -9.650 10.160 ;
        RECT -12.835 9.865 -11.605 9.960 ;
        RECT -8.890 9.695 -8.660 10.515 ;
        RECT -8.390 10.495 -8.160 10.710 ;
        RECT -8.490 9.865 -8.160 10.495 ;
        RECT -7.745 9.695 -7.455 10.420 ;
        RECT -28.070 9.525 -26.690 9.695 ;
        RECT -24.390 9.525 -23.010 9.695 ;
        RECT -20.250 9.525 -18.870 9.695 ;
        RECT -17.030 9.525 -15.650 9.695 ;
        RECT -13.350 9.525 -11.510 9.695 ;
        RECT -9.210 9.525 -7.370 9.695 ;
        RECT -25.880 8.555 -25.420 8.725 ;
        RECT -25.240 8.575 -23.860 8.745 ;
        RECT -21.390 8.625 -20.010 8.795 ;
        RECT -25.795 7.830 -25.505 8.555 ;
        RECT -25.155 7.775 -24.845 8.575 ;
        RECT -24.640 8.260 -23.945 8.405 ;
        RECT -24.640 8.060 -22.950 8.260 ;
        RECT -24.640 7.775 -23.945 8.060 ;
        RECT -21.305 7.825 -20.995 8.625 ;
        RECT -20.790 8.210 -20.095 8.455 ;
        RECT -20.790 8.010 -18.800 8.210 ;
        RECT -20.790 7.825 -20.095 8.010 ;
        RECT -25.145 7.560 -24.810 7.605 ;
        RECT -26.300 7.360 -24.810 7.560 ;
        RECT -25.145 7.335 -24.810 7.360 ;
        RECT -24.640 7.175 -24.470 7.775 ;
        RECT -21.295 7.610 -20.960 7.655 ;
        RECT -24.300 7.560 -23.965 7.585 ;
        RECT -24.300 7.360 -22.350 7.560 ;
        RECT -22.050 7.410 -20.960 7.610 ;
        RECT -21.295 7.385 -20.960 7.410 ;
        RECT -24.300 7.335 -23.965 7.360 ;
        RECT -25.795 6.005 -25.505 7.170 ;
        RECT -25.155 6.025 -24.875 7.165 ;
        RECT -24.705 6.195 -24.375 7.175 ;
        RECT -24.205 6.025 -23.945 7.165 ;
        RECT -23.275 7.060 -23.075 7.360 ;
        RECT -20.790 7.225 -20.620 7.825 ;
        RECT -20.450 7.595 -20.115 7.635 ;
        RECT -20.450 7.425 -19.515 7.595 ;
        RECT 10.995 7.525 11.165 12.045 ;
        RECT 12.720 10.700 14.500 10.870 ;
        RECT 12.720 8.880 12.890 10.700 ;
        RECT 13.445 10.190 13.775 10.360 ;
        RECT 13.290 9.560 13.460 10.020 ;
        RECT 13.760 9.560 13.930 10.020 ;
        RECT 13.445 9.220 13.775 9.390 ;
        RECT 14.330 8.880 14.500 10.700 ;
        RECT 12.720 8.710 14.500 8.880 ;
        RECT 16.065 7.525 16.235 12.045 ;
        RECT -20.450 7.385 -20.115 7.425 ;
        RECT 10.995 7.355 16.235 7.525 ;
        RECT 20.830 8.730 22.610 8.900 ;
        RECT -21.305 6.075 -21.025 7.215 ;
        RECT -20.855 6.245 -20.525 7.225 ;
        RECT -20.355 6.075 -20.095 7.215 ;
        RECT 20.830 6.700 21.000 8.730 ;
        RECT 21.555 8.220 21.885 8.390 ;
        RECT 21.400 7.425 21.570 8.005 ;
        RECT 21.870 7.425 22.040 8.005 ;
        RECT 21.555 7.040 21.885 7.210 ;
        RECT 22.440 6.700 22.610 8.730 ;
        RECT 138.630 7.035 139.720 7.145 ;
        RECT 138.295 6.865 140.045 7.035 ;
        RECT 157.780 6.865 158.630 6.925 ;
        RECT -14.610 6.435 -12.310 6.605 ;
        RECT -11.690 6.435 -11.230 6.605 ;
        RECT 20.830 6.530 22.610 6.700 ;
        RECT 120.400 6.695 121.260 6.815 ;
        RECT 119.945 6.525 121.695 6.695 ;
        RECT -25.880 5.835 -25.420 6.005 ;
        RECT -25.240 5.855 -23.860 6.025 ;
        RECT -21.390 5.905 -20.010 6.075 ;
        RECT -16.100 5.760 -15.900 6.410 ;
        RECT -16.100 5.560 -15.150 5.760 ;
        RECT -14.525 5.295 -14.265 6.435 ;
        RECT -14.095 5.465 -13.765 6.265 ;
        RECT -13.595 5.635 -13.425 6.435 ;
        RECT -13.225 5.465 -12.895 6.265 ;
        RECT -12.695 5.635 -12.415 6.435 ;
        RECT -14.095 5.295 -12.815 5.465 ;
        RECT -17.060 5.060 -14.940 5.070 ;
        RECT -14.500 5.060 -14.215 5.125 ;
        RECT -17.060 4.860 -14.200 5.060 ;
        RECT -17.060 4.850 -14.940 4.860 ;
        RECT -14.500 4.795 -14.215 4.860 ;
        RECT -14.015 4.795 -13.635 5.125 ;
        RECT -13.465 4.795 -13.155 5.125 ;
        RECT -16.000 4.210 -14.900 4.410 ;
        RECT -15.995 2.865 -15.805 4.210 ;
        RECT -14.520 3.885 -14.185 4.625 ;
        RECT -14.015 4.100 -13.800 4.795 ;
        RECT -13.465 4.625 -13.260 4.795 ;
        RECT -12.985 4.625 -12.815 5.295 ;
        RECT -12.635 5.060 -12.395 5.465 ;
        RECT -11.605 5.270 -11.315 6.435 ;
        RECT -12.635 4.860 -9.850 5.060 ;
        RECT -12.635 4.795 -12.395 4.860 ;
        RECT -13.610 4.100 -13.260 4.625 ;
        RECT -13.090 4.055 -12.395 4.625 ;
        RECT -11.605 3.885 -11.315 4.610 ;
        RECT 119.945 4.125 120.115 6.525 ;
        RECT 120.655 6.015 120.985 6.185 ;
        RECT 120.515 4.805 120.685 5.845 ;
        RECT 120.955 4.805 121.125 5.845 ;
        RECT 120.655 4.465 120.985 4.635 ;
        RECT 121.525 4.125 121.695 6.525 ;
        RECT 125.430 6.395 126.260 6.475 ;
        RECT 119.945 3.955 121.695 4.125 ;
        RECT 124.965 6.225 126.715 6.395 ;
        RECT -14.610 3.715 -12.310 3.885 ;
        RECT -11.690 3.715 -11.230 3.885 ;
        RECT 124.965 3.825 125.135 6.225 ;
        RECT 125.675 5.715 126.005 5.885 ;
        RECT 125.535 4.505 125.705 5.545 ;
        RECT 125.975 4.505 126.145 5.545 ;
        RECT 125.675 4.165 126.005 4.335 ;
        RECT 126.545 3.825 126.715 6.225 ;
        RECT 34.705 3.575 39.945 3.745 ;
        RECT 124.965 3.655 126.715 3.825 ;
        RECT 131.755 4.915 134.495 5.085 ;
        RECT 26.060 3.020 27.840 3.190 ;
        RECT 5.230 2.500 7.010 2.670 ;
        RECT 5.230 0.470 5.400 2.500 ;
        RECT 5.955 1.990 6.285 2.160 ;
        RECT 5.800 1.195 5.970 1.775 ;
        RECT 6.270 1.195 6.440 1.775 ;
        RECT 5.955 0.810 6.285 0.980 ;
        RECT 6.840 0.470 7.010 2.500 ;
        RECT 5.230 0.300 7.010 0.470 ;
        RECT 13.590 2.570 15.370 2.740 ;
        RECT 13.590 0.540 13.760 2.570 ;
        RECT 14.315 2.060 14.645 2.230 ;
        RECT 14.160 1.265 14.330 1.845 ;
        RECT 14.630 1.265 14.800 1.845 ;
        RECT 14.315 0.880 14.645 1.050 ;
        RECT 15.200 0.540 15.370 2.570 ;
        RECT 26.060 1.200 26.230 3.020 ;
        RECT 26.785 2.510 27.115 2.680 ;
        RECT 26.630 1.880 26.800 2.340 ;
        RECT 27.100 1.880 27.270 2.340 ;
        RECT 26.785 1.540 27.115 1.710 ;
        RECT 27.670 1.200 27.840 3.020 ;
        RECT 26.060 1.030 27.840 1.200 ;
        RECT 13.590 0.370 15.370 0.540 ;
        RECT -27.150 -0.675 -25.770 -0.505 ;
        RECT -23.470 -0.675 -22.090 -0.505 ;
        RECT -19.330 -0.675 -17.950 -0.505 ;
        RECT -16.110 -0.675 -14.730 -0.505 ;
        RECT -12.430 -0.675 -10.590 -0.505 ;
        RECT -8.290 -0.675 -6.910 -0.505 ;
        RECT -6.620 -0.665 -6.160 -0.495 ;
        RECT -26.810 -1.815 -26.600 -0.675 ;
        RECT -26.430 -1.825 -26.100 -0.845 ;
        RECT -23.385 -1.815 -23.105 -0.675 ;
        RECT -22.935 -1.825 -22.605 -0.845 ;
        RECT -22.435 -1.815 -22.175 -0.675 ;
        RECT -18.990 -1.815 -18.780 -0.675 ;
        RECT -18.610 -1.825 -18.280 -0.845 ;
        RECT -15.770 -1.815 -15.560 -0.675 ;
        RECT -15.390 -1.825 -15.060 -0.845 ;
        RECT -12.340 -1.815 -12.085 -0.675 ;
        RECT -11.915 -1.645 -11.585 -0.845 ;
        RECT -11.415 -1.475 -11.185 -0.675 ;
        RECT -11.015 -1.645 -10.685 -0.845 ;
        RECT -11.915 -1.815 -10.685 -1.645 ;
        RECT -7.950 -1.815 -7.740 -0.675 ;
        RECT -27.800 -1.995 -26.530 -1.990 ;
        RECT -27.800 -2.190 -26.500 -1.995 ;
        RECT -26.830 -2.235 -26.500 -2.190 ;
        RECT -26.330 -2.040 -26.100 -1.825 ;
        RECT -23.375 -2.040 -23.040 -1.985 ;
        RECT -26.330 -2.240 -23.040 -2.040 ;
        RECT -26.830 -3.225 -26.600 -2.405 ;
        RECT -26.330 -2.425 -26.100 -2.240 ;
        RECT -23.375 -2.255 -23.040 -2.240 ;
        RECT -22.870 -2.425 -22.700 -1.825 ;
        RECT -22.530 -1.990 -22.195 -1.985 ;
        RECT -18.510 -1.990 -18.280 -1.825 ;
        RECT -22.530 -2.190 -21.450 -1.990 ;
        RECT -19.850 -1.995 -18.750 -1.990 ;
        RECT -18.510 -1.995 -15.550 -1.990 ;
        RECT -19.850 -2.190 -18.680 -1.995 ;
        RECT -22.530 -2.235 -22.195 -2.190 ;
        RECT -26.430 -3.055 -26.100 -2.425 ;
        RECT -23.385 -3.225 -23.075 -2.425 ;
        RECT -22.870 -2.690 -22.175 -2.425 ;
        RECT -20.500 -2.690 -20.300 -2.240 ;
        RECT -19.850 -2.690 -19.650 -2.190 ;
        RECT -19.010 -2.235 -18.680 -2.190 ;
        RECT -18.510 -2.190 -15.460 -1.995 ;
        RECT -22.870 -2.890 -19.650 -2.690 ;
        RECT -22.870 -3.055 -22.175 -2.890 ;
        RECT -19.010 -3.225 -18.780 -2.405 ;
        RECT -18.510 -2.425 -18.280 -2.190 ;
        RECT -15.790 -2.235 -15.460 -2.190 ;
        RECT -15.290 -2.040 -15.060 -1.825 ;
        RECT -12.320 -2.040 -12.100 -1.985 ;
        RECT -15.290 -2.240 -13.200 -2.040 ;
        RECT -13.000 -2.240 -12.100 -2.040 ;
        RECT -18.610 -3.055 -18.280 -2.425 ;
        RECT -15.790 -3.225 -15.560 -2.405 ;
        RECT -15.290 -2.425 -15.060 -2.240 ;
        RECT -15.390 -3.055 -15.060 -2.425 ;
        RECT -12.320 -2.565 -12.100 -2.240 ;
        RECT -11.915 -2.715 -11.735 -1.815 ;
        RECT -7.570 -1.825 -7.240 -0.845 ;
        RECT -11.565 -2.545 -11.190 -1.985 ;
        RECT -10.985 -2.055 -10.675 -1.985 ;
        RECT -9.200 -2.055 -8.350 -2.040 ;
        RECT -7.970 -2.055 -7.640 -1.995 ;
        RECT -10.985 -2.225 -9.920 -2.055 ;
        RECT -9.200 -2.225 -7.640 -2.055 ;
        RECT -10.985 -2.315 -10.675 -2.225 ;
        RECT -9.200 -2.240 -8.350 -2.225 ;
        RECT -7.970 -2.235 -7.640 -2.225 ;
        RECT -7.470 -2.040 -7.240 -1.825 ;
        RECT -6.535 -1.830 -6.245 -0.665 ;
        RECT 5.120 -0.980 6.900 -0.810 ;
        RECT -11.015 -2.715 -10.685 -2.485 ;
        RECT -12.340 -3.225 -12.085 -2.735 ;
        RECT -11.915 -2.740 -10.685 -2.715 ;
        RECT -8.550 -2.740 -8.350 -2.240 ;
        RECT -7.470 -2.240 -4.800 -2.040 ;
        RECT -11.915 -2.940 -8.350 -2.740 ;
        RECT -11.915 -3.055 -10.685 -2.940 ;
        RECT -7.970 -3.225 -7.740 -2.405 ;
        RECT -7.470 -2.425 -7.240 -2.240 ;
        RECT -7.570 -3.055 -7.240 -2.425 ;
        RECT -6.535 -3.215 -6.245 -2.490 ;
        RECT 5.120 -2.800 5.290 -0.980 ;
        RECT 5.845 -1.490 6.175 -1.320 ;
        RECT 5.690 -2.120 5.860 -1.660 ;
        RECT 6.160 -2.120 6.330 -1.660 ;
        RECT 5.845 -2.460 6.175 -2.290 ;
        RECT 6.730 -2.800 6.900 -0.980 ;
        RECT 34.705 -0.945 34.875 3.575 ;
        RECT 36.460 2.240 38.240 2.410 ;
        RECT 36.460 0.420 36.630 2.240 ;
        RECT 37.185 1.730 37.515 1.900 ;
        RECT 37.030 1.100 37.200 1.560 ;
        RECT 37.500 1.100 37.670 1.560 ;
        RECT 37.185 0.760 37.515 0.930 ;
        RECT 38.070 0.420 38.240 2.240 ;
        RECT 36.460 0.250 38.240 0.420 ;
        RECT 39.775 -0.945 39.945 3.575 ;
        RECT 131.755 3.505 131.925 4.915 ;
        RECT 134.325 4.635 134.495 4.915 ;
        RECT 132.265 4.045 132.435 4.375 ;
        RECT 132.605 4.345 133.645 4.515 ;
        RECT 132.605 3.905 133.645 4.075 ;
        RECT 133.815 4.045 133.985 4.375 ;
        RECT 134.325 3.665 134.555 4.635 ;
        RECT 138.295 4.465 138.465 6.865 ;
        RECT 139.005 6.355 139.335 6.525 ;
        RECT 138.865 5.145 139.035 6.185 ;
        RECT 139.305 5.145 139.475 6.185 ;
        RECT 139.005 4.805 139.335 4.975 ;
        RECT 139.875 4.465 140.045 6.865 ;
        RECT 144.215 6.655 145.085 6.725 ;
        RECT 157.330 6.695 159.080 6.865 ;
        RECT 138.295 4.295 140.045 4.465 ;
        RECT 143.775 6.485 145.525 6.655 ;
        RECT 143.775 4.085 143.945 6.485 ;
        RECT 144.485 5.975 144.815 6.145 ;
        RECT 144.345 4.765 144.515 5.805 ;
        RECT 144.785 4.765 144.955 5.805 ;
        RECT 144.485 4.425 144.815 4.595 ;
        RECT 145.355 4.085 145.525 6.485 ;
        RECT 143.775 3.915 145.525 4.085 ;
        RECT 151.555 5.495 154.295 5.665 ;
        RECT 151.555 4.085 151.725 5.495 ;
        RECT 154.125 5.185 154.295 5.495 ;
        RECT 152.065 4.625 152.235 4.955 ;
        RECT 152.405 4.925 153.445 5.095 ;
        RECT 152.405 4.485 153.445 4.655 ;
        RECT 153.615 4.625 153.785 4.955 ;
        RECT 154.125 4.325 154.380 5.185 ;
        RECT 154.125 4.085 154.295 4.325 ;
        RECT 157.330 4.295 157.500 6.695 ;
        RECT 158.040 6.185 158.370 6.355 ;
        RECT 157.900 4.975 158.070 6.015 ;
        RECT 158.340 4.975 158.510 6.015 ;
        RECT 158.040 4.635 158.370 4.805 ;
        RECT 158.910 4.295 159.080 6.695 ;
        RECT 157.330 4.125 159.080 4.295 ;
        RECT 151.555 3.915 154.295 4.085 ;
        RECT 134.325 3.505 134.495 3.665 ;
        RECT 131.755 3.335 134.495 3.505 ;
        RECT 119.975 3.135 121.725 3.305 ;
        RECT 57.670 -0.835 58.660 -0.695 ;
        RECT 65.260 -0.785 66.250 -0.645 ;
        RECT 72.870 -0.765 73.860 -0.625 ;
        RECT 23.375 -1.225 28.615 -1.055 ;
        RECT 34.705 -1.115 39.945 -0.945 ;
        RECT 57.290 -1.005 59.070 -0.835 ;
        RECT 5.120 -2.970 6.900 -2.800 ;
        RECT 12.055 -2.535 17.295 -2.365 ;
        RECT -27.150 -3.395 -25.770 -3.225 ;
        RECT -23.470 -3.395 -22.090 -3.225 ;
        RECT -19.330 -3.395 -17.950 -3.225 ;
        RECT -16.110 -3.395 -14.730 -3.225 ;
        RECT -12.430 -3.395 -10.590 -3.225 ;
        RECT -8.290 -3.395 -6.910 -3.225 ;
        RECT -6.620 -3.385 -6.160 -3.215 ;
        RECT -23.930 -3.785 -22.550 -3.615 ;
        RECT -23.845 -4.340 -23.150 -3.955 ;
        RECT -24.900 -4.540 -23.150 -4.340 ;
        RECT -23.845 -4.585 -23.150 -4.540 ;
        RECT -22.945 -4.585 -22.635 -3.785 ;
        RECT -20.700 -3.845 -19.320 -3.675 ;
        RECT -20.615 -4.190 -19.920 -4.015 ;
        RECT -22.350 -4.390 -19.920 -4.190 ;
        RECT -23.825 -4.855 -23.490 -4.775 ;
        RECT -25.135 -5.025 -23.490 -4.855 ;
        RECT -23.320 -5.185 -23.150 -4.585 ;
        RECT -22.980 -4.790 -22.645 -4.755 ;
        RECT -22.350 -4.790 -22.150 -4.390 ;
        RECT -22.980 -4.990 -22.150 -4.790 ;
        RECT -22.980 -5.025 -22.645 -4.990 ;
        RECT -23.845 -6.335 -23.585 -5.195 ;
        RECT -23.415 -6.165 -23.085 -5.185 ;
        RECT -22.915 -6.335 -22.635 -5.195 ;
        RECT -21.800 -5.690 -21.600 -4.390 ;
        RECT -20.615 -4.645 -19.920 -4.390 ;
        RECT -19.715 -4.645 -19.405 -3.845 ;
        RECT -19.110 -3.915 -18.650 -3.745 ;
        RECT -19.025 -4.640 -18.735 -3.915 ;
        RECT -20.595 -4.855 -20.260 -4.835 ;
        RECT -21.135 -5.025 -20.260 -4.855 ;
        RECT -20.595 -5.085 -20.260 -5.025 ;
        RECT -20.090 -5.245 -19.920 -4.645 ;
        RECT -19.750 -4.840 -19.415 -4.815 ;
        RECT -19.750 -5.040 -18.000 -4.840 ;
        RECT -19.750 -5.085 -19.415 -5.040 ;
        RECT -23.930 -6.505 -22.550 -6.335 ;
        RECT -20.615 -6.395 -20.355 -5.255 ;
        RECT -20.185 -6.225 -19.855 -5.245 ;
        RECT -19.685 -6.395 -19.405 -5.255 ;
        RECT -20.700 -6.565 -19.320 -6.395 ;
        RECT -19.025 -6.465 -18.735 -5.300 ;
        RECT -19.110 -6.635 -18.650 -6.465 ;
        RECT 12.055 -7.055 12.225 -2.535 ;
        RECT 13.700 -3.900 15.480 -3.730 ;
        RECT 13.700 -5.720 13.870 -3.900 ;
        RECT 14.425 -4.410 14.755 -4.240 ;
        RECT 14.270 -5.040 14.440 -4.580 ;
        RECT 14.740 -5.040 14.910 -4.580 ;
        RECT 14.425 -5.380 14.755 -5.210 ;
        RECT 15.310 -5.720 15.480 -3.900 ;
        RECT 13.700 -5.890 15.480 -5.720 ;
        RECT 17.125 -7.055 17.295 -2.535 ;
        RECT 23.375 -5.745 23.545 -1.225 ;
        RECT 25.160 -2.590 26.940 -2.420 ;
        RECT 25.160 -4.410 25.330 -2.590 ;
        RECT 25.885 -3.100 26.215 -2.930 ;
        RECT 25.730 -3.730 25.900 -3.270 ;
        RECT 26.200 -3.730 26.370 -3.270 ;
        RECT 25.885 -4.070 26.215 -3.900 ;
        RECT 26.770 -4.410 26.940 -2.590 ;
        RECT 25.160 -4.580 26.940 -4.410 ;
        RECT 28.445 -5.745 28.615 -1.225 ;
        RECT 23.375 -5.915 28.615 -5.745 ;
        RECT 48.530 -2.755 50.310 -2.585 ;
        RECT 48.530 -6.045 48.700 -2.755 ;
        RECT 49.255 -3.265 49.585 -3.095 ;
        RECT 49.100 -5.320 49.270 -3.480 ;
        RECT 49.570 -5.320 49.740 -3.480 ;
        RECT 49.255 -5.705 49.585 -5.535 ;
        RECT 50.140 -6.045 50.310 -2.755 ;
        RECT 57.290 -3.215 57.460 -1.005 ;
        RECT 58.015 -1.515 58.345 -1.345 ;
        RECT 57.860 -2.490 58.030 -1.730 ;
        RECT 58.330 -2.490 58.500 -1.730 ;
        RECT 58.015 -2.875 58.345 -2.705 ;
        RECT 58.900 -3.215 59.070 -1.005 ;
        RECT 57.290 -3.385 59.070 -3.215 ;
        RECT 64.880 -0.955 66.660 -0.785 ;
        RECT 64.880 -3.165 65.050 -0.955 ;
        RECT 65.605 -1.465 65.935 -1.295 ;
        RECT 65.450 -2.440 65.620 -1.680 ;
        RECT 65.920 -2.440 66.090 -1.680 ;
        RECT 65.605 -2.825 65.935 -2.655 ;
        RECT 66.490 -3.165 66.660 -0.955 ;
        RECT 64.880 -3.335 66.660 -3.165 ;
        RECT 72.490 -0.935 74.270 -0.765 ;
        RECT 80.870 -0.805 81.860 -0.665 ;
        RECT 88.680 -0.785 89.670 -0.645 ;
        RECT 72.490 -3.145 72.660 -0.935 ;
        RECT 73.215 -1.445 73.545 -1.275 ;
        RECT 73.060 -2.420 73.230 -1.660 ;
        RECT 73.530 -2.420 73.700 -1.660 ;
        RECT 73.215 -2.805 73.545 -2.635 ;
        RECT 74.100 -3.145 74.270 -0.935 ;
        RECT 72.490 -3.315 74.270 -3.145 ;
        RECT 80.490 -0.975 82.270 -0.805 ;
        RECT 80.490 -3.185 80.660 -0.975 ;
        RECT 81.215 -1.485 81.545 -1.315 ;
        RECT 81.060 -2.460 81.230 -1.700 ;
        RECT 81.530 -2.460 81.700 -1.700 ;
        RECT 81.215 -2.845 81.545 -2.675 ;
        RECT 82.100 -3.185 82.270 -0.975 ;
        RECT 80.490 -3.355 82.270 -3.185 ;
        RECT 88.300 -0.955 90.080 -0.785 ;
        RECT 96.270 -0.805 97.260 -0.665 ;
        RECT 88.300 -3.165 88.470 -0.955 ;
        RECT 89.025 -1.465 89.355 -1.295 ;
        RECT 88.870 -2.440 89.040 -1.680 ;
        RECT 89.340 -2.440 89.510 -1.680 ;
        RECT 89.025 -2.825 89.355 -2.655 ;
        RECT 89.910 -3.165 90.080 -0.955 ;
        RECT 88.300 -3.335 90.080 -3.165 ;
        RECT 95.890 -0.975 97.670 -0.805 ;
        RECT 103.660 -0.835 104.650 -0.695 ;
        RECT 95.890 -3.185 96.060 -0.975 ;
        RECT 96.615 -1.485 96.945 -1.315 ;
        RECT 96.460 -2.460 96.630 -1.700 ;
        RECT 96.930 -2.460 97.100 -1.700 ;
        RECT 96.615 -2.845 96.945 -2.675 ;
        RECT 97.500 -3.185 97.670 -0.975 ;
        RECT 95.890 -3.355 97.670 -3.185 ;
        RECT 103.280 -1.005 105.060 -0.835 ;
        RECT 103.280 -3.215 103.450 -1.005 ;
        RECT 104.005 -1.515 104.335 -1.345 ;
        RECT 103.850 -2.490 104.020 -1.730 ;
        RECT 104.320 -2.490 104.490 -1.730 ;
        RECT 104.005 -2.875 104.335 -2.705 ;
        RECT 104.890 -3.215 105.060 -1.005 ;
        RECT 119.975 -0.855 120.145 3.135 ;
        RECT 120.685 2.625 121.015 2.795 ;
        RECT 120.545 -0.130 120.715 2.410 ;
        RECT 120.985 -0.130 121.155 2.410 ;
        RECT 120.685 -0.515 121.015 -0.345 ;
        RECT 121.555 -0.855 121.725 3.135 ;
        RECT 138.355 3.275 140.105 3.445 ;
        RECT 119.975 -1.025 121.725 -0.855 ;
        RECT 124.995 2.905 126.745 3.075 ;
        RECT 120.350 -1.175 121.320 -1.025 ;
        RECT 124.995 -1.085 125.165 2.905 ;
        RECT 125.705 2.395 126.035 2.565 ;
        RECT 125.565 -0.360 125.735 2.180 ;
        RECT 126.005 -0.360 126.175 2.180 ;
        RECT 125.705 -0.745 126.035 -0.575 ;
        RECT 125.415 -1.085 126.325 -1.075 ;
        RECT 126.575 -1.085 126.745 2.905 ;
        RECT 131.005 2.155 135.335 2.325 ;
        RECT 131.005 1.995 131.175 2.155 ;
        RECT 130.895 0.885 131.175 1.995 ;
        RECT 131.515 1.285 131.685 1.615 ;
        RECT 131.900 1.585 134.440 1.755 ;
        RECT 131.900 1.145 134.440 1.315 ;
        RECT 134.655 1.285 134.825 1.615 ;
        RECT 131.005 0.745 131.175 0.885 ;
        RECT 135.165 0.745 135.335 2.155 ;
        RECT 131.005 0.575 135.335 0.745 ;
        RECT 138.355 -0.715 138.525 3.275 ;
        RECT 139.065 2.765 139.395 2.935 ;
        RECT 138.925 0.010 139.095 2.550 ;
        RECT 139.365 0.010 139.535 2.550 ;
        RECT 139.065 -0.375 139.395 -0.205 ;
        RECT 139.935 -0.715 140.105 3.275 ;
        RECT 138.355 -0.885 140.105 -0.715 ;
        RECT 143.805 3.265 145.555 3.435 ;
        RECT 143.805 -0.725 143.975 3.265 ;
        RECT 144.515 2.755 144.845 2.925 ;
        RECT 144.375 0.000 144.545 2.540 ;
        RECT 144.815 0.000 144.985 2.540 ;
        RECT 144.515 -0.385 144.845 -0.215 ;
        RECT 145.385 -0.725 145.555 3.265 ;
        RECT 157.310 3.065 159.060 3.235 ;
        RECT 150.705 2.635 155.035 2.805 ;
        RECT 150.705 2.335 150.875 2.635 ;
        RECT 150.640 1.485 150.875 2.335 ;
        RECT 151.215 1.765 151.385 2.095 ;
        RECT 151.600 2.065 154.140 2.235 ;
        RECT 151.600 1.625 154.140 1.795 ;
        RECT 154.355 1.765 154.525 2.095 ;
        RECT 150.705 1.225 150.875 1.485 ;
        RECT 154.865 1.225 155.035 2.635 ;
        RECT 150.705 1.055 155.035 1.225 ;
        RECT 138.805 -1.025 139.775 -0.885 ;
        RECT 143.805 -0.895 145.555 -0.725 ;
        RECT 144.195 -0.935 145.135 -0.895 ;
        RECT 157.310 -0.925 157.480 3.065 ;
        RECT 158.020 2.555 158.350 2.725 ;
        RECT 157.880 -0.200 158.050 2.340 ;
        RECT 158.320 -0.200 158.490 2.340 ;
        RECT 158.020 -0.585 158.350 -0.415 ;
        RECT 158.890 -0.925 159.060 3.065 ;
        RECT 124.995 -1.255 126.745 -1.085 ;
        RECT 157.310 -1.095 159.060 -0.925 ;
        RECT 157.680 -1.225 158.650 -1.095 ;
        RECT 125.415 -1.415 126.325 -1.255 ;
        RECT 110.290 -2.965 111.130 -2.885 ;
        RECT 103.280 -3.385 105.060 -3.215 ;
        RECT 109.800 -3.135 111.580 -2.965 ;
        RECT 48.530 -6.215 50.310 -6.045 ;
        RECT 57.290 -3.825 59.070 -3.655 ;
        RECT 57.290 -6.035 57.460 -3.825 ;
        RECT 58.015 -4.335 58.345 -4.165 ;
        RECT 57.860 -5.310 58.030 -4.550 ;
        RECT 58.330 -5.310 58.500 -4.550 ;
        RECT 58.015 -5.695 58.345 -5.525 ;
        RECT 58.900 -6.035 59.070 -3.825 ;
        RECT 57.290 -6.205 59.070 -6.035 ;
        RECT 64.880 -3.775 66.660 -3.605 ;
        RECT 64.880 -5.985 65.050 -3.775 ;
        RECT 65.605 -4.285 65.935 -4.115 ;
        RECT 65.450 -5.260 65.620 -4.500 ;
        RECT 65.920 -5.260 66.090 -4.500 ;
        RECT 65.605 -5.645 65.935 -5.475 ;
        RECT 66.490 -5.985 66.660 -3.775 ;
        RECT 64.880 -6.155 66.660 -5.985 ;
        RECT 72.490 -3.755 74.270 -3.585 ;
        RECT 72.490 -5.965 72.660 -3.755 ;
        RECT 73.215 -4.265 73.545 -4.095 ;
        RECT 73.060 -5.240 73.230 -4.480 ;
        RECT 73.530 -5.240 73.700 -4.480 ;
        RECT 73.215 -5.625 73.545 -5.455 ;
        RECT 74.100 -5.965 74.270 -3.755 ;
        RECT 72.490 -6.135 74.270 -5.965 ;
        RECT 80.490 -3.795 82.270 -3.625 ;
        RECT 80.490 -6.005 80.660 -3.795 ;
        RECT 81.215 -4.305 81.545 -4.135 ;
        RECT 81.060 -5.280 81.230 -4.520 ;
        RECT 81.530 -5.280 81.700 -4.520 ;
        RECT 81.215 -5.665 81.545 -5.495 ;
        RECT 82.100 -6.005 82.270 -3.795 ;
        RECT 80.490 -6.175 82.270 -6.005 ;
        RECT 88.300 -3.775 90.080 -3.605 ;
        RECT 88.300 -5.985 88.470 -3.775 ;
        RECT 89.025 -4.285 89.355 -4.115 ;
        RECT 88.870 -5.260 89.040 -4.500 ;
        RECT 89.340 -5.260 89.510 -4.500 ;
        RECT 89.025 -5.645 89.355 -5.475 ;
        RECT 89.910 -5.985 90.080 -3.775 ;
        RECT 88.300 -6.155 90.080 -5.985 ;
        RECT 95.890 -3.795 97.670 -3.625 ;
        RECT 95.890 -6.005 96.060 -3.795 ;
        RECT 96.615 -4.305 96.945 -4.135 ;
        RECT 96.460 -5.280 96.630 -4.520 ;
        RECT 96.930 -5.280 97.100 -4.520 ;
        RECT 96.615 -5.665 96.945 -5.495 ;
        RECT 97.500 -6.005 97.670 -3.795 ;
        RECT 95.890 -6.175 97.670 -6.005 ;
        RECT 103.280 -3.825 105.060 -3.655 ;
        RECT 103.280 -6.035 103.450 -3.825 ;
        RECT 104.005 -4.335 104.335 -4.165 ;
        RECT 103.850 -5.310 104.020 -4.550 ;
        RECT 104.320 -5.310 104.490 -4.550 ;
        RECT 104.005 -5.695 104.335 -5.525 ;
        RECT 104.890 -6.035 105.060 -3.825 ;
        RECT 109.800 -5.345 109.970 -3.135 ;
        RECT 110.525 -3.645 110.855 -3.475 ;
        RECT 110.370 -4.620 110.540 -3.860 ;
        RECT 110.840 -4.620 111.010 -3.860 ;
        RECT 110.525 -5.005 110.855 -4.835 ;
        RECT 111.410 -5.345 111.580 -3.135 ;
        RECT 109.800 -5.515 111.580 -5.345 ;
        RECT 121.965 -4.685 124.705 -4.515 ;
        RECT 103.280 -6.205 105.060 -6.035 ;
        RECT 121.965 -6.095 122.135 -4.685 ;
        RECT 124.535 -4.995 124.705 -4.685 ;
        RECT 122.475 -5.555 122.645 -5.225 ;
        RECT 122.815 -5.255 123.855 -5.085 ;
        RECT 122.815 -5.695 123.855 -5.525 ;
        RECT 124.025 -5.555 124.195 -5.225 ;
        RECT 124.515 -5.875 124.715 -4.995 ;
        RECT 142.155 -5.435 144.895 -5.265 ;
        RECT 124.535 -6.095 124.705 -5.875 ;
        RECT 121.965 -6.265 124.705 -6.095 ;
        RECT 109.750 -6.525 111.530 -6.355 ;
        RECT 12.055 -7.225 17.295 -7.055 ;
        RECT 57.300 -6.975 59.080 -6.805 ;
        RECT 48.520 -7.615 50.300 -7.445 ;
        RECT 48.520 -9.435 48.690 -7.615 ;
        RECT 49.245 -8.125 49.575 -7.955 ;
        RECT 49.090 -8.755 49.260 -8.295 ;
        RECT 49.560 -8.755 49.730 -8.295 ;
        RECT 49.245 -9.095 49.575 -8.925 ;
        RECT 50.130 -9.435 50.300 -7.615 ;
        RECT 57.300 -8.795 57.470 -6.975 ;
        RECT 58.025 -7.485 58.355 -7.315 ;
        RECT 57.870 -8.115 58.040 -7.655 ;
        RECT 58.340 -8.115 58.510 -7.655 ;
        RECT 58.025 -8.455 58.355 -8.285 ;
        RECT 58.910 -8.795 59.080 -6.975 ;
        RECT 57.300 -8.965 59.080 -8.795 ;
        RECT 64.890 -6.925 66.670 -6.755 ;
        RECT 64.890 -8.745 65.060 -6.925 ;
        RECT 65.615 -7.435 65.945 -7.265 ;
        RECT 65.460 -8.065 65.630 -7.605 ;
        RECT 65.930 -8.065 66.100 -7.605 ;
        RECT 65.615 -8.405 65.945 -8.235 ;
        RECT 66.500 -8.745 66.670 -6.925 ;
        RECT 64.890 -8.915 66.670 -8.745 ;
        RECT 72.500 -6.905 74.280 -6.735 ;
        RECT 72.500 -8.725 72.670 -6.905 ;
        RECT 73.225 -7.415 73.555 -7.245 ;
        RECT 73.070 -8.045 73.240 -7.585 ;
        RECT 73.540 -8.045 73.710 -7.585 ;
        RECT 73.225 -8.385 73.555 -8.215 ;
        RECT 74.110 -8.725 74.280 -6.905 ;
        RECT 72.500 -8.895 74.280 -8.725 ;
        RECT 80.500 -6.945 82.280 -6.775 ;
        RECT 80.500 -8.765 80.670 -6.945 ;
        RECT 81.225 -7.455 81.555 -7.285 ;
        RECT 81.070 -8.085 81.240 -7.625 ;
        RECT 81.540 -8.085 81.710 -7.625 ;
        RECT 81.225 -8.425 81.555 -8.255 ;
        RECT 82.110 -8.765 82.280 -6.945 ;
        RECT 80.500 -8.935 82.280 -8.765 ;
        RECT 88.310 -6.925 90.090 -6.755 ;
        RECT 88.310 -8.745 88.480 -6.925 ;
        RECT 89.035 -7.435 89.365 -7.265 ;
        RECT 88.880 -8.065 89.050 -7.605 ;
        RECT 89.350 -8.065 89.520 -7.605 ;
        RECT 89.035 -8.405 89.365 -8.235 ;
        RECT 89.920 -8.745 90.090 -6.925 ;
        RECT 88.310 -8.915 90.090 -8.745 ;
        RECT 95.900 -6.945 97.680 -6.775 ;
        RECT 95.900 -8.765 96.070 -6.945 ;
        RECT 96.625 -7.455 96.955 -7.285 ;
        RECT 96.470 -8.085 96.640 -7.625 ;
        RECT 96.940 -8.085 97.110 -7.625 ;
        RECT 96.625 -8.425 96.955 -8.255 ;
        RECT 97.510 -8.765 97.680 -6.945 ;
        RECT 95.900 -8.935 97.680 -8.765 ;
        RECT 103.290 -6.975 105.070 -6.805 ;
        RECT 103.290 -8.795 103.460 -6.975 ;
        RECT 104.015 -7.485 104.345 -7.315 ;
        RECT 103.860 -8.115 104.030 -7.655 ;
        RECT 104.330 -8.115 104.500 -7.655 ;
        RECT 104.015 -8.455 104.345 -8.285 ;
        RECT 104.900 -8.795 105.070 -6.975 ;
        RECT 109.750 -8.345 109.920 -6.525 ;
        RECT 110.475 -7.035 110.805 -6.865 ;
        RECT 110.320 -7.665 110.490 -7.205 ;
        RECT 110.790 -7.665 110.960 -7.205 ;
        RECT 110.475 -8.005 110.805 -7.835 ;
        RECT 111.360 -8.345 111.530 -6.525 ;
        RECT 142.155 -6.845 142.325 -5.435 ;
        RECT 144.725 -5.705 144.895 -5.435 ;
        RECT 142.665 -6.305 142.835 -5.975 ;
        RECT 143.005 -6.005 144.045 -5.835 ;
        RECT 143.005 -6.445 144.045 -6.275 ;
        RECT 144.215 -6.305 144.385 -5.975 ;
        RECT 144.725 -6.605 145.095 -5.705 ;
        RECT 144.725 -6.845 144.895 -6.605 ;
        RECT 142.155 -7.015 144.895 -6.845 ;
        RECT 109.750 -8.515 111.530 -8.345 ;
        RECT 121.045 -7.555 125.375 -7.385 ;
        RECT 110.140 -8.625 111.150 -8.515 ;
        RECT 103.290 -8.965 105.070 -8.795 ;
        RECT 121.045 -8.965 121.215 -7.555 ;
        RECT 121.555 -8.425 121.725 -8.095 ;
        RECT 121.940 -8.125 124.480 -7.955 ;
        RECT 121.940 -8.565 124.480 -8.395 ;
        RECT 124.695 -8.425 124.865 -8.095 ;
        RECT 125.205 -8.965 125.375 -7.555 ;
        RECT 141.395 -8.275 145.725 -8.105 ;
        RECT 141.395 -8.615 141.565 -8.275 ;
        RECT 121.045 -9.135 125.375 -8.965 ;
        RECT 48.520 -9.605 50.300 -9.435 ;
        RECT 57.310 -9.405 59.090 -9.235 ;
        RECT 17.190 -10.800 33.930 -10.630 ;
        RECT 17.190 -12.240 17.360 -10.800 ;
        RECT 17.700 -11.685 17.870 -11.355 ;
        RECT 18.040 -11.370 33.080 -11.200 ;
        RECT 18.040 -11.840 33.080 -11.670 ;
        RECT 33.250 -11.685 33.420 -11.355 ;
        RECT 33.760 -12.240 33.930 -10.800 ;
        RECT 57.310 -11.225 57.480 -9.405 ;
        RECT 58.035 -9.915 58.365 -9.745 ;
        RECT 57.880 -10.545 58.050 -10.085 ;
        RECT 58.350 -10.545 58.520 -10.085 ;
        RECT 58.035 -10.885 58.365 -10.715 ;
        RECT 57.740 -11.225 58.690 -11.205 ;
        RECT 58.920 -11.225 59.090 -9.405 ;
        RECT 57.310 -11.395 59.090 -11.225 ;
        RECT 64.900 -9.355 66.680 -9.185 ;
        RECT 64.900 -11.175 65.070 -9.355 ;
        RECT 65.625 -9.865 65.955 -9.695 ;
        RECT 65.470 -10.495 65.640 -10.035 ;
        RECT 65.940 -10.495 66.110 -10.035 ;
        RECT 65.625 -10.835 65.955 -10.665 ;
        RECT 65.330 -11.175 66.280 -11.155 ;
        RECT 66.510 -11.175 66.680 -9.355 ;
        RECT 64.900 -11.345 66.680 -11.175 ;
        RECT 72.510 -9.335 74.290 -9.165 ;
        RECT 72.510 -11.155 72.680 -9.335 ;
        RECT 73.235 -9.845 73.565 -9.675 ;
        RECT 73.080 -10.475 73.250 -10.015 ;
        RECT 73.550 -10.475 73.720 -10.015 ;
        RECT 73.235 -10.815 73.565 -10.645 ;
        RECT 72.940 -11.155 73.890 -11.135 ;
        RECT 74.120 -11.155 74.290 -9.335 ;
        RECT 72.510 -11.325 74.290 -11.155 ;
        RECT 80.510 -9.375 82.290 -9.205 ;
        RECT 80.510 -11.195 80.680 -9.375 ;
        RECT 81.235 -9.885 81.565 -9.715 ;
        RECT 81.080 -10.515 81.250 -10.055 ;
        RECT 81.550 -10.515 81.720 -10.055 ;
        RECT 81.235 -10.855 81.565 -10.685 ;
        RECT 80.940 -11.195 81.890 -11.175 ;
        RECT 82.120 -11.195 82.290 -9.375 ;
        RECT 80.510 -11.365 82.290 -11.195 ;
        RECT 88.320 -9.355 90.100 -9.185 ;
        RECT 88.320 -11.175 88.490 -9.355 ;
        RECT 89.045 -9.865 89.375 -9.695 ;
        RECT 88.890 -10.495 89.060 -10.035 ;
        RECT 89.360 -10.495 89.530 -10.035 ;
        RECT 89.045 -10.835 89.375 -10.665 ;
        RECT 88.750 -11.175 89.700 -11.155 ;
        RECT 89.930 -11.175 90.100 -9.355 ;
        RECT 88.320 -11.345 90.100 -11.175 ;
        RECT 95.910 -9.375 97.690 -9.205 ;
        RECT 95.910 -11.195 96.080 -9.375 ;
        RECT 96.635 -9.885 96.965 -9.715 ;
        RECT 96.480 -10.515 96.650 -10.055 ;
        RECT 96.950 -10.515 97.120 -10.055 ;
        RECT 96.635 -10.855 96.965 -10.685 ;
        RECT 96.340 -11.195 97.290 -11.175 ;
        RECT 97.520 -11.195 97.690 -9.375 ;
        RECT 95.910 -11.365 97.690 -11.195 ;
        RECT 103.300 -9.405 105.080 -9.235 ;
        RECT 141.255 -9.365 141.565 -8.615 ;
        RECT 141.905 -9.145 142.075 -8.815 ;
        RECT 142.290 -8.845 144.830 -8.675 ;
        RECT 142.290 -9.285 144.830 -9.115 ;
        RECT 145.045 -9.145 145.215 -8.815 ;
        RECT 103.300 -11.225 103.470 -9.405 ;
        RECT 104.025 -9.915 104.355 -9.745 ;
        RECT 103.870 -10.545 104.040 -10.085 ;
        RECT 104.340 -10.545 104.510 -10.085 ;
        RECT 104.025 -10.885 104.355 -10.715 ;
        RECT 103.730 -11.225 104.680 -11.205 ;
        RECT 104.910 -11.225 105.080 -9.405 ;
        RECT 141.395 -9.685 141.565 -9.365 ;
        RECT 145.555 -9.685 145.725 -8.275 ;
        RECT 141.395 -9.855 145.725 -9.685 ;
        RECT 103.300 -11.395 105.080 -11.225 ;
        RECT 17.190 -12.410 33.930 -12.240 ;
      LAYER met1 ;
        RECT 77.790 86.440 88.560 86.880 ;
        RECT 71.750 75.600 76.560 76.120 ;
        RECT 71.750 61.320 72.270 75.600 ;
        RECT 71.720 60.320 76.460 61.320 ;
        RECT 71.750 55.180 72.270 60.320 ;
        RECT 71.720 54.660 72.300 55.180 ;
        RECT 64.660 52.330 65.180 52.360 ;
        RECT 64.660 51.810 75.880 52.330 ;
        RECT 64.660 51.780 65.180 51.810 ;
        RECT 71.750 35.900 72.270 50.870 ;
        RECT 67.370 35.380 72.270 35.900 ;
        RECT 75.360 33.870 75.880 51.810 ;
        RECT 60.670 33.350 75.880 33.870 ;
        RECT 60.670 32.150 61.190 33.350 ;
        RECT 60.710 31.250 61.030 32.150 ;
        RECT 60.680 29.145 61.060 31.250 ;
        RECT 60.680 25.340 61.060 27.445 ;
        RECT 60.710 24.290 61.030 25.340 ;
        RECT 60.710 23.940 61.010 24.290 ;
        RECT 60.670 23.500 61.010 23.940 ;
        RECT 42.230 23.165 42.460 23.210 ;
        RECT 42.230 22.935 44.905 23.165 ;
        RECT 42.230 21.870 42.460 22.935 ;
        RECT 44.675 22.470 44.905 22.935 ;
        RECT 60.710 23.100 61.010 23.500 ;
        RECT -2.070 20.320 -1.790 21.700 ;
        RECT 25.260 21.640 43.330 21.870 ;
        RECT -1.500 21.170 16.570 21.400 ;
        RECT 15.220 20.520 15.480 21.170 ;
        RECT 16.980 20.320 17.140 20.340 ;
        RECT 43.590 20.320 43.870 21.670 ;
        RECT 44.090 20.650 45.100 22.470 ;
        RECT -2.070 20.040 43.870 20.320 ;
        RECT 15.190 19.470 16.780 19.730 ;
        RECT 11.960 18.140 12.960 18.530 ;
        RECT -0.640 17.790 12.960 18.140 ;
        RECT 16.980 18.010 17.140 20.040 ;
        RECT 17.770 19.730 18.030 19.760 ;
        RECT 17.770 19.470 29.030 19.730 ;
        RECT 17.770 19.440 18.030 19.470 ;
        RECT 22.330 18.615 22.660 18.630 ;
        RECT 22.330 18.285 25.925 18.615 ;
        RECT -0.640 15.755 -0.290 17.790 ;
        RECT 11.960 17.420 12.960 17.790 ;
        RECT 16.900 17.750 17.220 18.010 ;
        RECT 22.330 17.680 22.660 18.285 ;
        RECT 22.160 17.420 22.660 17.680 ;
        RECT 4.510 17.390 22.660 17.420 ;
        RECT 4.510 16.870 22.740 17.390 ;
        RECT 3.750 16.490 4.070 16.520 ;
        RECT 4.600 16.490 6.460 16.870 ;
        RECT 3.750 16.300 6.460 16.490 ;
        RECT 3.750 16.290 6.240 16.300 ;
        RECT 3.750 16.260 4.070 16.290 ;
        RECT 4.680 16.270 6.240 16.290 ;
        RECT 11.430 16.040 11.710 16.870 ;
        RECT 22.345 16.765 22.740 16.870 ;
        RECT 24.770 16.765 25.090 16.790 ;
        RECT 22.345 16.555 25.090 16.765 ;
        RECT 16.930 16.140 17.190 16.460 ;
        RECT 23.305 16.300 23.515 16.555 ;
        RECT 24.770 16.530 25.090 16.555 ;
        RECT 26.805 16.390 27.035 19.470 ;
        RECT 28.850 16.970 29.030 19.470 ;
        RECT 44.535 19.325 44.865 20.650 ;
        RECT 36.865 18.995 55.615 19.325 ;
        RECT 29.645 18.615 29.975 18.645 ;
        RECT 36.865 18.615 37.195 18.995 ;
        RECT 29.645 18.285 37.195 18.615 ;
        RECT 29.645 18.255 29.975 18.285 ;
        RECT 60.710 18.140 61.030 23.100 ;
        RECT 39.820 17.820 61.030 18.140 ;
        RECT 28.850 16.790 29.720 16.970 ;
        RECT 28.850 16.600 29.030 16.790 ;
        RECT -8.345 15.405 -0.290 15.755 ;
        RECT -22.580 14.560 -22.320 14.620 ;
        RECT -10.360 14.560 -10.040 14.590 ;
        RECT -22.580 14.360 -10.040 14.560 ;
        RECT -22.580 14.300 -22.320 14.360 ;
        RECT -10.360 14.330 -10.040 14.360 ;
        RECT -18.140 13.250 -17.140 14.110 ;
        RECT -8.345 13.250 -7.995 15.405 ;
        RECT -1.250 13.680 -0.930 13.710 ;
        RECT -1.900 13.480 -0.930 13.680 ;
        RECT -27.800 12.770 -7.660 13.250 ;
        RECT -27.800 12.570 -7.100 12.770 ;
        RECT -28.070 12.430 -7.100 12.570 ;
        RECT -28.070 12.090 -26.690 12.430 ;
        RECT -24.390 12.090 -23.010 12.430 ;
        RECT -20.250 12.090 -18.870 12.430 ;
        RECT -17.030 12.090 -15.650 12.430 ;
        RECT -13.350 12.090 -11.510 12.430 ;
        RECT -22.610 11.630 -22.290 11.890 ;
        RECT -10.330 11.850 -10.070 12.170 ;
        RECT -9.210 12.090 -7.370 12.430 ;
        RECT -14.860 11.810 -14.540 11.840 ;
        RECT -30.450 10.980 -29.450 11.390 ;
        RECT -31.700 10.910 -29.450 10.980 ;
        RECT -28.780 10.910 -28.520 10.970 ;
        RECT -22.550 10.925 -22.350 11.630 ;
        RECT -21.550 11.110 -21.250 11.790 ;
        RECT -14.860 11.610 -12.250 11.810 ;
        RECT -14.860 11.580 -14.540 11.610 ;
        RECT -31.700 10.730 -28.520 10.910 ;
        RECT -30.450 10.710 -28.520 10.730 ;
        RECT -30.450 10.390 -29.450 10.710 ;
        RECT -28.780 10.650 -28.520 10.710 ;
        RECT -22.595 10.695 -22.305 10.925 ;
        RECT -21.580 10.810 -21.220 11.110 ;
        RECT -12.450 10.855 -12.250 11.610 ;
        RECT -10.300 11.520 -10.100 11.850 ;
        RECT -10.330 11.200 -10.070 11.520 ;
        RECT -7.030 10.910 -6.770 10.970 ;
        RECT -1.900 10.910 -1.700 13.480 ;
        RECT -1.250 13.450 -0.930 13.480 ;
        RECT -12.465 10.565 -12.235 10.855 ;
        RECT -7.030 10.710 -1.700 10.910 ;
        RECT -10.875 10.640 -10.615 10.675 ;
        RECT -7.030 10.650 -6.770 10.710 ;
        RECT -10.905 10.385 -10.590 10.640 ;
        RECT -10.875 10.355 -10.615 10.385 ;
        RECT -15.060 10.010 -14.740 10.040 ;
        RECT -13.995 10.010 -13.705 10.025 ;
        RECT -28.070 9.510 -26.690 9.850 ;
        RECT -24.390 9.510 -23.010 9.850 ;
        RECT -20.250 9.510 -18.870 9.850 ;
        RECT -17.030 9.510 -15.650 9.850 ;
        RECT -15.060 9.810 -13.705 10.010 ;
        RECT -15.060 9.780 -14.740 9.810 ;
        RECT -13.995 9.795 -13.705 9.810 ;
        RECT -13.350 9.510 -11.510 9.850 ;
        RECT -9.210 9.510 -7.370 9.850 ;
        RECT -28.070 9.370 -7.370 9.510 ;
        RECT -27.800 9.030 -7.100 9.370 ;
        RECT -27.800 8.690 -7.660 9.030 ;
        RECT -25.880 8.400 -25.420 8.690 ;
        RECT -25.240 8.420 -23.860 8.690 ;
        RECT -21.390 8.470 -20.010 8.690 ;
        RECT -23.180 8.000 -22.920 8.320 ;
        RECT -22.580 8.000 -22.320 8.320 ;
        RECT -19.760 8.180 -19.440 8.440 ;
        RECT -22.550 7.620 -22.350 8.000 ;
        RECT -26.345 7.345 -26.055 7.575 ;
        RECT -26.300 4.460 -26.100 7.345 ;
        RECT -23.290 7.290 -23.030 7.320 ;
        RECT -22.580 7.300 -22.320 7.620 ;
        RECT -22.080 7.350 -21.820 7.670 ;
        RECT -19.680 7.655 -19.520 8.180 ;
        RECT -19.030 7.950 -18.770 8.270 ;
        RECT -17.680 8.010 -16.680 8.690 ;
        RECT -15.060 8.180 -14.740 8.440 ;
        RECT -19.715 7.365 -19.485 7.655 ;
        RECT -23.320 7.030 -23.030 7.290 ;
        RECT -23.290 7.000 -23.030 7.030 ;
        RECT -23.255 6.355 -22.935 6.395 ;
        RECT -22.040 6.355 -21.855 7.350 ;
        RECT -25.880 5.970 -25.420 6.160 ;
        RECT -25.240 5.970 -23.860 6.180 ;
        RECT -23.255 6.170 -21.855 6.355 ;
        RECT -23.255 6.135 -22.935 6.170 ;
        RECT -21.390 5.970 -20.010 6.230 ;
        RECT -25.880 5.680 -19.520 5.970 ;
        RECT -25.500 5.290 -19.520 5.680 ;
        RECT -22.280 4.610 -21.280 5.290 ;
        RECT -19.000 4.460 -18.800 7.950 ;
        RECT -15.000 7.860 -14.800 8.180 ;
        RECT -15.000 7.660 -9.850 7.860 ;
        RECT -16.130 7.000 -15.870 7.320 ;
        RECT -16.100 6.455 -15.900 7.000 ;
        RECT -13.900 6.760 -12.900 7.510 ;
        RECT -16.115 6.165 -15.885 6.455 ;
        RECT -14.610 6.280 -11.230 6.760 ;
        RECT -12.450 6.260 -11.480 6.280 ;
        RECT -15.380 5.760 -15.120 5.820 ;
        RECT -15.380 5.560 -13.750 5.760 ;
        RECT -15.380 5.500 -15.120 5.560 ;
        RECT -13.950 5.105 -13.750 5.560 ;
        RECT -10.050 5.105 -9.850 7.660 ;
        RECT -17.095 4.845 -16.805 5.075 ;
        RECT -26.300 4.260 -18.800 4.460 ;
        RECT -23.250 3.735 -22.930 3.995 ;
        RECT -23.180 2.465 -22.995 3.735 ;
        RECT -21.060 3.220 -20.740 3.240 ;
        RECT -17.060 3.220 -16.840 4.845 ;
        RECT -13.965 4.815 -13.735 5.105 ;
        RECT -10.065 4.815 -9.835 5.105 ;
        RECT -12.990 4.510 -12.700 4.535 ;
        RECT -12.275 4.510 -12.015 4.575 ;
        RECT -15.130 4.410 -14.870 4.470 ;
        RECT -13.595 4.410 -13.305 4.425 ;
        RECT -15.130 4.210 -13.305 4.410 ;
        RECT -12.990 4.325 -12.015 4.510 ;
        RECT -12.990 4.305 -12.700 4.325 ;
        RECT -12.275 4.255 -12.015 4.325 ;
        RECT -15.130 4.150 -14.870 4.210 ;
        RECT -13.595 4.195 -13.305 4.210 ;
        RECT -12.450 4.040 -11.480 4.060 ;
        RECT -14.610 3.560 -11.230 4.040 ;
        RECT -0.640 3.785 -0.290 15.405 ;
        RECT 2.730 15.770 5.640 16.000 ;
        RECT 11.410 15.780 13.750 16.040 ;
        RECT 2.730 14.795 2.960 15.770 ;
        RECT 5.315 15.760 5.605 15.770 ;
        RECT 11.410 15.680 11.710 15.780 ;
        RECT 3.750 15.410 4.070 15.440 ;
        RECT 5.110 15.410 5.340 15.555 ;
        RECT 3.750 15.210 5.340 15.410 ;
        RECT 3.750 15.180 4.070 15.210 ;
        RECT 5.110 15.015 5.340 15.210 ;
        RECT 5.580 15.380 5.810 15.555 ;
        RECT 5.580 15.160 6.850 15.380 ;
        RECT 5.580 15.015 5.810 15.160 ;
        RECT 5.315 14.795 5.605 14.810 ;
        RECT 2.730 14.580 5.605 14.795 ;
        RECT 2.730 14.565 5.595 14.580 ;
        RECT 0.680 13.910 1.680 14.280 ;
        RECT 2.730 13.910 2.960 14.565 ;
        RECT 0.030 13.680 0.290 13.740 ;
        RECT 0.680 13.690 2.960 13.910 ;
        RECT 0.680 13.680 1.680 13.690 ;
        RECT 0.030 13.480 1.680 13.680 ;
        RECT 0.030 13.420 0.290 13.480 ;
        RECT 0.680 13.280 1.680 13.480 ;
        RECT 2.170 6.620 2.390 13.690 ;
        RECT 2.730 13.085 2.960 13.690 ;
        RECT 4.210 13.920 4.530 13.940 ;
        RECT 6.630 13.920 6.850 15.160 ;
        RECT 11.410 14.580 11.670 15.680 ;
        RECT 13.240 15.420 13.470 15.605 ;
        RECT 12.200 15.260 13.470 15.420 ;
        RECT 12.200 14.010 12.360 15.260 ;
        RECT 13.240 15.065 13.470 15.260 ;
        RECT 13.710 15.480 13.940 15.605 ;
        RECT 13.710 15.270 15.100 15.480 ;
        RECT 13.710 15.065 13.940 15.270 ;
        RECT 12.600 14.870 12.860 14.900 ;
        RECT 12.600 14.610 13.760 14.870 ;
        RECT 12.600 14.580 12.860 14.610 ;
        RECT 12.810 14.250 14.370 14.350 ;
        RECT 12.610 14.060 14.500 14.250 ;
        RECT 12.610 14.010 14.650 14.060 ;
        RECT 4.210 13.700 9.950 13.920 ;
        RECT 12.200 13.850 14.650 14.010 ;
        RECT 14.330 13.800 14.650 13.850 ;
        RECT 4.210 13.680 4.530 13.700 ;
        RECT 2.730 12.855 5.635 13.085 ;
        RECT 9.730 12.900 9.950 13.700 ;
        RECT 14.890 12.945 15.100 15.270 ;
        RECT 15.550 13.770 15.810 14.090 ;
        RECT 11.465 12.900 15.100 12.945 ;
        RECT 2.730 12.065 2.960 12.855 ;
        RECT 5.335 12.820 5.625 12.855 ;
        RECT 9.730 12.735 15.100 12.900 ;
        RECT 15.600 13.100 15.760 13.770 ;
        RECT 16.980 13.100 17.140 16.140 ;
        RECT 23.120 16.070 24.680 16.300 ;
        RECT 26.790 16.070 27.050 16.390 ;
        RECT 28.810 16.280 29.070 16.600 ;
        RECT 29.540 16.430 29.720 16.790 ;
        RECT 29.410 16.420 30.330 16.430 ;
        RECT 29.410 16.220 30.390 16.420 ;
        RECT 29.695 16.190 30.390 16.220 ;
        RECT 23.750 15.570 25.650 15.820 ;
        RECT 23.755 15.560 24.045 15.570 ;
        RECT 23.550 15.140 23.780 15.355 ;
        RECT 15.600 12.940 17.140 13.100 ;
        RECT 22.450 14.940 23.780 15.140 ;
        RECT 9.730 12.680 11.675 12.735 ;
        RECT 4.210 12.530 4.530 12.550 ;
        RECT 5.130 12.530 5.360 12.660 ;
        RECT 4.210 12.310 5.360 12.530 ;
        RECT 4.210 12.290 4.530 12.310 ;
        RECT 5.130 12.240 5.360 12.310 ;
        RECT 5.600 12.630 5.830 12.660 ;
        RECT 5.600 12.380 6.880 12.630 ;
        RECT 5.600 12.240 5.830 12.380 ;
        RECT 5.335 12.065 5.625 12.080 ;
        RECT 2.730 11.835 5.635 12.065 ;
        RECT 6.630 11.615 6.880 12.380 ;
        RECT 5.715 11.570 6.880 11.615 ;
        RECT 4.620 11.365 6.880 11.570 ;
        RECT 4.620 10.900 6.480 11.365 ;
        RECT 4.650 6.620 4.970 6.640 ;
        RECT 2.170 6.400 4.970 6.620 ;
        RECT 4.650 6.380 4.970 6.400 ;
        RECT 5.350 5.170 5.630 10.900 ;
        RECT 10.810 10.420 11.090 10.450 ;
        RECT 9.960 10.140 11.090 10.420 ;
        RECT 9.960 9.440 10.240 10.140 ;
        RECT 10.810 10.110 11.090 10.140 ;
        RECT 11.465 9.865 11.675 12.680 ;
        RECT 11.900 10.140 13.790 10.420 ;
        RECT 13.260 9.865 13.490 10.000 ;
        RECT 11.465 9.655 13.490 9.865 ;
        RECT 13.260 9.580 13.490 9.655 ;
        RECT 13.730 9.810 13.960 10.000 ;
        RECT 15.600 9.810 15.760 12.940 ;
        RECT 22.450 12.390 22.650 14.940 ;
        RECT 23.550 14.815 23.780 14.940 ;
        RECT 24.020 15.190 24.250 15.355 ;
        RECT 25.400 15.245 25.650 15.570 ;
        RECT 27.660 15.690 29.780 15.930 ;
        RECT 27.660 15.245 27.900 15.690 ;
        RECT 29.465 15.680 29.755 15.690 ;
        RECT 24.770 15.190 25.090 15.215 ;
        RECT 24.020 14.980 25.090 15.190 ;
        RECT 24.020 14.815 24.250 14.980 ;
        RECT 24.770 14.955 25.090 14.980 ;
        RECT 25.400 14.995 27.900 15.245 ;
        RECT 28.780 15.270 29.100 15.310 ;
        RECT 29.260 15.270 29.490 15.475 ;
        RECT 28.780 15.090 29.490 15.270 ;
        RECT 28.780 15.050 29.100 15.090 ;
        RECT 25.400 14.700 25.650 14.995 ;
        RECT 27.660 14.740 27.900 14.995 ;
        RECT 29.260 14.935 29.490 15.090 ;
        RECT 29.730 15.340 29.960 15.475 ;
        RECT 29.730 15.130 31.320 15.340 ;
        RECT 29.730 14.935 29.960 15.130 ;
        RECT 27.660 14.730 29.750 14.740 ;
        RECT 25.400 14.665 25.680 14.700 ;
        RECT 23.765 14.610 25.680 14.665 ;
        RECT 23.755 14.415 25.680 14.610 ;
        RECT 27.660 14.500 29.755 14.730 ;
        RECT 23.755 14.380 24.045 14.415 ;
        RECT 25.480 12.390 25.680 14.415 ;
        RECT 26.790 14.160 27.050 14.480 ;
        RECT 13.730 9.650 15.760 9.810 ;
        RECT 18.030 12.190 25.680 12.390 ;
        RECT 13.730 9.580 13.960 9.650 ;
        RECT 9.960 9.160 13.800 9.440 ;
        RECT 6.180 6.620 6.440 6.670 ;
        RECT 8.990 6.620 9.310 6.640 ;
        RECT 6.180 6.400 9.310 6.620 ;
        RECT 6.180 6.350 6.440 6.400 ;
        RECT 8.990 6.380 9.310 6.400 ;
        RECT 9.960 5.170 10.240 9.160 ;
        RECT 12.830 8.890 14.390 8.910 ;
        RECT 14.900 8.890 15.060 9.650 ;
        RECT 12.830 8.730 15.060 8.890 ;
        RECT 12.830 8.680 14.390 8.730 ;
        RECT 18.030 7.490 18.230 12.190 ;
        RECT 19.130 8.420 21.850 8.430 ;
        RECT 19.130 8.210 21.865 8.420 ;
        RECT 18.000 7.170 18.260 7.490 ;
        RECT 19.130 7.190 19.350 8.210 ;
        RECT 21.575 8.190 21.865 8.210 ;
        RECT 21.370 7.880 21.600 7.985 ;
        RECT 21.840 7.880 22.070 7.985 ;
        RECT 22.410 7.880 22.640 8.790 ;
        RECT 26.805 7.880 27.035 14.160 ;
        RECT 31.110 9.440 31.320 15.130 ;
        RECT 39.820 9.440 40.140 17.820 ;
        RECT 55.225 16.375 55.615 16.705 ;
        RECT 55.255 16.000 55.585 16.375 ;
        RECT 55.190 14.760 61.570 16.000 ;
        RECT 55.255 13.265 55.585 14.760 ;
        RECT 77.790 12.540 78.230 86.440 ;
        RECT 80.920 60.290 81.920 61.350 ;
        RECT 43.640 12.100 78.230 12.540 ;
        RECT 81.200 12.230 81.640 60.290 ;
        RECT 91.620 38.120 140.735 38.390 ;
        RECT 91.620 25.830 91.890 38.120 ;
        RECT 103.095 36.535 106.595 36.605 ;
        RECT 103.095 36.335 133.165 36.535 ;
        RECT 103.095 29.805 103.365 36.335 ;
        RECT 106.220 36.265 133.165 36.335 ;
        RECT 106.085 32.260 106.395 32.690 ;
        RECT 107.760 32.260 108.020 32.320 ;
        RECT 104.635 32.060 108.020 32.260 ;
        RECT 126.185 32.210 127.185 33.240 ;
        RECT 104.635 30.430 104.835 32.060 ;
        RECT 106.085 32.050 106.395 32.060 ;
        RECT 107.760 32.000 108.020 32.060 ;
        RECT 126.475 31.785 126.795 32.210 ;
        RECT 106.845 31.510 110.165 31.710 ;
        RECT 106.845 30.620 107.045 31.510 ;
        RECT 108.315 30.820 108.905 31.130 ;
        RECT 104.635 30.140 104.865 30.430 ;
        RECT 105.070 30.390 107.570 30.620 ;
        RECT 107.760 30.520 108.020 30.820 ;
        RECT 104.635 30.130 104.835 30.140 ;
        RECT 105.070 29.950 107.570 30.180 ;
        RECT 107.725 30.090 108.055 30.520 ;
        RECT 94.045 29.535 103.365 29.805 ;
        RECT 91.160 25.350 92.160 25.830 ;
        RECT 87.090 25.010 92.160 25.350 ;
        RECT 85.470 18.655 86.470 19.020 ;
        RECT 84.005 18.365 86.470 18.655 ;
        RECT 43.640 9.440 44.080 12.100 ;
        RECT 81.200 11.790 83.270 12.230 ;
        RECT 81.200 10.680 81.640 11.790 ;
        RECT 50.410 10.240 81.640 10.680 ;
        RECT 48.070 9.440 49.070 9.650 ;
        RECT 31.080 9.080 49.070 9.440 ;
        RECT 21.370 7.650 27.035 7.880 ;
        RECT 21.370 7.445 21.600 7.650 ;
        RECT 21.840 7.445 22.070 7.650 ;
        RECT 21.575 7.190 21.865 7.240 ;
        RECT 19.110 6.970 21.890 7.190 ;
        RECT 10.840 6.620 11.100 6.670 ;
        RECT 19.110 6.620 19.330 6.970 ;
        RECT 22.410 6.640 22.640 7.650 ;
        RECT 10.840 6.400 19.330 6.620 ;
        RECT 10.840 6.350 11.100 6.400 ;
        RECT 17.970 5.500 18.290 5.760 ;
        RECT 18.030 5.170 18.230 5.500 ;
        RECT 5.320 5.125 18.390 5.170 ;
        RECT 1.165 4.815 18.390 5.125 ;
        RECT -21.060 3.000 -16.840 3.220 ;
        RECT -16.045 3.055 -15.755 3.075 ;
        RECT -14.060 3.055 -13.740 3.090 ;
        RECT -21.060 2.980 -20.740 3.000 ;
        RECT -16.045 2.865 -13.740 3.055 ;
        RECT -16.045 2.845 -15.755 2.865 ;
        RECT -14.060 2.830 -13.740 2.865 ;
        RECT -13.350 2.760 -12.350 3.560 ;
        RECT -0.670 3.435 -0.260 3.785 ;
        RECT -11.560 2.465 -11.240 2.505 ;
        RECT -23.180 2.280 -11.240 2.465 ;
        RECT -23.180 0.605 -22.995 2.280 ;
        RECT -11.560 2.245 -11.240 2.280 ;
        RECT -29.040 0.420 -22.995 0.605 ;
        RECT -21.650 1.410 -9.000 1.610 ;
        RECT -21.650 0.520 -21.450 1.410 ;
        RECT -31.450 -1.990 -30.450 -1.690 ;
        RECT -29.880 -1.990 -29.620 -1.930 ;
        RECT -31.450 -2.190 -29.620 -1.990 ;
        RECT -31.450 -2.690 -30.450 -2.190 ;
        RECT -29.880 -2.250 -29.620 -2.190 ;
        RECT -31.175 -10.535 -30.845 -2.690 ;
        RECT -29.035 -6.560 -28.865 0.420 ;
        RECT -21.680 0.200 -21.420 0.520 ;
        RECT -16.760 -0.015 -15.760 0.850 ;
        RECT -9.200 0.540 -9.000 1.410 ;
        RECT -9.260 0.280 -8.940 0.540 ;
        RECT -26.870 -0.150 -6.730 -0.015 ;
        RECT -26.870 -0.340 -6.180 -0.150 ;
        RECT -26.870 -0.350 -6.160 -0.340 ;
        RECT -27.150 -0.820 -6.160 -0.350 ;
        RECT -27.150 -0.830 -6.550 -0.820 ;
        RECT -26.870 -0.835 -6.550 -0.830 ;
        RECT -6.800 -0.840 -6.550 -0.835 ;
        RECT -21.710 -1.320 -21.390 -1.060 ;
        RECT -13.450 -1.240 -11.250 -1.040 ;
        RECT -28.510 -1.990 -28.190 -1.960 ;
        RECT -27.830 -1.990 -27.570 -1.930 ;
        RECT -21.650 -1.975 -21.450 -1.320 ;
        RECT -20.530 -1.570 -20.270 -1.250 ;
        RECT -21.060 -1.790 -20.740 -1.760 ;
        RECT -20.500 -1.790 -20.300 -1.570 ;
        RECT -28.510 -2.190 -27.570 -1.990 ;
        RECT -28.510 -2.220 -28.190 -2.190 ;
        RECT -27.830 -2.250 -27.570 -2.190 ;
        RECT -21.695 -2.205 -21.405 -1.975 ;
        RECT -21.060 -1.990 -20.300 -1.790 ;
        RECT -21.060 -2.020 -20.740 -1.990 ;
        RECT -20.500 -2.225 -20.300 -1.990 ;
        RECT -13.450 -2.010 -13.250 -1.240 ;
        RECT -20.545 -2.455 -20.255 -2.225 ;
        RECT -13.510 -2.270 -13.190 -2.010 ;
        RECT -13.045 -2.255 -12.755 -2.025 ;
        RECT -11.450 -2.045 -11.250 -1.240 ;
        RECT -10.165 -1.320 -9.845 -1.060 ;
        RECT -9.230 -1.300 -8.970 -0.980 ;
        RECT -10.090 -1.995 -9.920 -1.320 ;
        RECT -9.200 -1.980 -9.000 -1.300 ;
        RECT -13.000 -2.610 -12.800 -2.255 ;
        RECT -11.465 -2.335 -11.235 -2.045 ;
        RECT -10.120 -2.285 -9.890 -1.995 ;
        RECT -9.230 -2.300 -8.970 -1.980 ;
        RECT -5.030 -2.040 -4.770 -1.980 ;
        RECT 0.470 -2.040 0.790 -2.010 ;
        RECT -5.030 -2.240 0.790 -2.040 ;
        RECT -5.030 -2.300 -4.770 -2.240 ;
        RECT 0.470 -2.270 0.790 -2.240 ;
        RECT -13.060 -2.870 -12.740 -2.610 ;
        RECT -6.800 -3.060 -6.500 -3.040 ;
        RECT -6.800 -3.070 -6.160 -3.060 ;
        RECT -27.150 -3.210 -6.160 -3.070 ;
        RECT -27.340 -3.525 -6.160 -3.210 ;
        RECT 1.165 -3.525 1.475 4.815 ;
        RECT 5.320 4.650 18.390 4.815 ;
        RECT 2.385 4.305 2.735 4.335 ;
        RECT 10.130 4.305 11.130 4.440 ;
        RECT 2.385 3.955 11.130 4.305 ;
        RECT 2.385 3.925 2.735 3.955 ;
        RECT 10.130 3.430 11.130 3.955 ;
        RECT 19.205 3.525 29.645 3.755 ;
        RECT 5.470 3.280 18.330 3.430 ;
        RECT 5.350 3.275 18.330 3.280 ;
        RECT 19.205 3.275 19.435 3.525 ;
        RECT 5.350 3.260 19.435 3.275 ;
        RECT 4.850 3.060 19.435 3.260 ;
        RECT 4.850 2.690 5.050 3.060 ;
        RECT 5.350 3.045 19.435 3.060 ;
        RECT 5.350 3.000 18.330 3.045 ;
        RECT 5.350 2.700 7.230 3.000 ;
        RECT 4.790 2.430 5.110 2.690 ;
        RECT 5.340 2.530 7.230 2.700 ;
        RECT 5.340 2.470 6.900 2.530 ;
        RECT 5.975 2.180 6.265 2.190 ;
        RECT 3.750 1.970 6.280 2.180 ;
        RECT 11.500 2.100 11.780 3.000 ;
        RECT 29.415 2.815 29.645 3.525 ;
        RECT 26.845 2.710 30.055 2.815 ;
        RECT 26.805 2.585 30.055 2.710 ;
        RECT 26.805 2.480 27.095 2.585 ;
        RECT 12.100 2.100 14.640 2.260 ;
        RECT 26.600 2.220 26.830 2.320 ;
        RECT 11.500 1.980 14.640 2.100 ;
        RECT 25.590 2.040 26.830 2.220 ;
        RECT 3.750 0.935 3.960 1.970 ;
        RECT 5.975 1.960 6.265 1.970 ;
        RECT 11.500 1.820 12.380 1.980 ;
        RECT 4.790 1.560 5.110 1.590 ;
        RECT 5.770 1.560 6.000 1.755 ;
        RECT 4.790 1.360 6.000 1.560 ;
        RECT 4.790 1.330 5.110 1.360 ;
        RECT 5.770 1.215 6.000 1.360 ;
        RECT 6.240 1.560 6.470 1.755 ;
        RECT 6.240 1.370 7.580 1.560 ;
        RECT 6.240 1.215 6.470 1.370 ;
        RECT 5.975 0.935 6.265 1.010 ;
        RECT 3.750 0.725 6.305 0.935 ;
        RECT 1.870 0.020 2.870 0.220 ;
        RECT 3.750 0.020 3.960 0.725 ;
        RECT 1.870 -0.260 3.960 0.020 ;
        RECT 7.390 0.180 7.580 1.370 ;
        RECT 12.100 0.780 12.380 1.820 ;
        RECT 14.130 1.570 14.360 1.825 ;
        RECT 12.950 1.390 14.360 1.570 ;
        RECT 12.950 0.230 13.130 1.390 ;
        RECT 14.130 1.285 14.360 1.390 ;
        RECT 14.600 1.670 14.830 1.825 ;
        RECT 14.600 1.500 16.160 1.670 ;
        RECT 14.600 1.285 14.830 1.500 ;
        RECT 13.290 1.090 13.570 1.120 ;
        RECT 13.290 0.810 14.710 1.090 ;
        RECT 13.290 0.780 13.570 0.810 ;
        RECT 13.700 0.420 15.260 0.570 ;
        RECT 13.530 0.400 15.370 0.420 ;
        RECT 13.530 0.270 15.470 0.400 ;
        RECT 13.530 0.230 15.730 0.270 ;
        RECT 7.390 -0.100 11.510 0.180 ;
        RECT 12.950 0.050 15.730 0.230 ;
        RECT 7.390 -0.255 7.580 -0.100 ;
        RECT 1.870 -0.780 2.870 -0.260 ;
        RECT 1.830 -2.040 2.090 -1.980 ;
        RECT 2.350 -2.040 2.550 -0.780 ;
        RECT 1.830 -2.240 2.550 -2.040 ;
        RECT 1.830 -2.300 2.090 -2.240 ;
        RECT -27.340 -3.835 1.475 -3.525 ;
        RECT -27.340 -3.890 -6.690 -3.835 ;
        RECT -23.930 -3.940 -22.550 -3.890 ;
        RECT -20.700 -4.000 -19.320 -3.890 ;
        RECT -19.110 -4.070 -18.650 -3.890 ;
        RECT -24.930 -4.600 -24.670 -4.280 ;
        RECT -21.210 -4.470 -20.890 -4.210 ;
        RECT -18.230 -4.400 -17.970 -4.080 ;
        RECT -21.135 -4.795 -20.965 -4.470 ;
        RECT -25.195 -5.055 -24.905 -4.825 ;
        RECT -25.130 -6.560 -24.970 -5.055 ;
        RECT -21.165 -5.085 -20.935 -4.795 ;
        RECT -18.200 -4.810 -18.000 -4.400 ;
        RECT -14.030 -4.450 -13.770 -4.130 ;
        RECT -18.260 -5.070 -17.940 -4.810 ;
        RECT -21.860 -5.490 -21.540 -5.460 ;
        RECT -14.000 -5.490 -13.800 -4.450 ;
        RECT -13.030 -4.550 -12.770 -4.230 ;
        RECT -9.700 -4.390 -8.700 -3.890 ;
        RECT -13.000 -5.490 -12.800 -4.550 ;
        RECT -21.860 -5.690 -12.800 -5.490 ;
        RECT -21.860 -5.720 -21.540 -5.690 ;
        RECT -29.035 -6.720 -24.970 -6.560 ;
        RECT -23.930 -6.610 -22.550 -6.180 ;
        RECT -20.700 -6.610 -19.320 -6.240 ;
        RECT -19.110 -6.610 -18.650 -6.310 ;
        RECT -29.035 -6.725 -28.865 -6.720 ;
        RECT -24.120 -6.790 -18.650 -6.610 ;
        RECT -24.120 -6.950 -19.060 -6.790 ;
        RECT -21.360 -7.870 -20.360 -6.950 ;
        RECT 1.165 -8.110 1.475 -3.835 ;
        RECT 3.140 -6.840 3.420 -0.260 ;
        RECT 3.750 -1.325 3.960 -0.260 ;
        RECT 5.045 -0.445 7.580 -0.255 ;
        RECT 5.045 -0.650 5.235 -0.445 ;
        RECT 5.010 -0.970 5.270 -0.650 ;
        RECT 5.865 -1.325 6.155 -1.290 ;
        RECT 3.750 -1.535 6.205 -1.325 ;
        RECT 11.230 -1.335 11.510 -0.100 ;
        RECT 15.380 0.010 15.730 0.050 ;
        RECT 15.380 -0.900 15.560 0.010 ;
        RECT 15.340 -1.220 15.600 -0.900 ;
        RECT 11.230 -1.385 13.140 -1.335 ;
        RECT 15.990 -1.385 16.160 1.500 ;
        RECT 25.590 1.190 25.770 2.040 ;
        RECT 26.600 1.900 26.830 2.040 ;
        RECT 27.070 2.260 27.300 2.320 ;
        RECT 28.350 2.260 28.560 2.585 ;
        RECT 27.070 2.050 28.560 2.260 ;
        RECT 27.070 1.900 27.300 2.050 ;
        RECT 26.805 1.710 27.095 1.740 ;
        RECT 27.490 1.710 28.455 1.765 ;
        RECT 26.805 1.535 28.455 1.710 ;
        RECT 26.805 1.510 27.095 1.535 ;
        RECT 28.225 1.425 28.455 1.535 ;
        RECT 29.825 1.425 30.055 2.585 ;
        RECT 31.110 2.715 31.320 9.080 ;
        RECT 48.070 8.630 49.070 9.080 ;
        RECT 48.550 6.120 48.890 8.630 ;
        RECT 44.390 5.780 48.890 6.120 ;
        RECT 50.410 5.490 50.850 10.240 ;
        RECT 40.950 5.050 50.850 5.490 ;
        RECT 51.405 8.925 55.615 9.255 ;
        RECT 35.900 2.715 36.220 2.740 ;
        RECT 31.110 2.505 36.220 2.715 ;
        RECT 35.900 2.480 36.220 2.505 ;
        RECT 32.800 1.710 37.570 1.940 ;
        RECT 32.800 1.425 33.030 1.710 ;
        RECT 37.205 1.700 37.495 1.710 ;
        RECT 26.170 1.190 27.730 1.230 ;
        RECT 28.225 1.195 33.030 1.425 ;
        RECT 20.240 1.010 27.730 1.190 ;
        RECT 20.240 0.730 20.420 1.010 ;
        RECT 26.170 1.000 27.730 1.010 ;
        RECT 32.800 0.915 33.030 1.195 ;
        RECT 35.900 1.425 36.220 1.450 ;
        RECT 37.000 1.425 37.230 1.540 ;
        RECT 35.900 1.215 37.230 1.425 ;
        RECT 35.900 1.190 36.220 1.215 ;
        RECT 37.000 1.120 37.230 1.215 ;
        RECT 37.470 1.485 37.700 1.540 ;
        RECT 37.470 1.295 38.645 1.485 ;
        RECT 37.470 1.120 37.700 1.295 ;
        RECT 37.205 0.915 37.495 0.960 ;
        RECT 20.200 0.410 20.460 0.730 ;
        RECT 32.800 0.685 37.565 0.915 ;
        RECT 36.570 0.405 38.130 0.450 ;
        RECT 38.455 0.405 38.645 1.295 ;
        RECT 16.390 0.230 16.650 0.300 ;
        RECT 16.390 0.050 22.340 0.230 ;
        RECT 36.570 0.220 38.645 0.405 ;
        RECT 16.390 -0.020 16.650 0.050 ;
        RECT 20.170 -0.620 20.490 -0.360 ;
        RECT 11.230 -1.500 16.160 -1.385 ;
        RECT 3.750 -2.315 3.960 -1.535 ;
        RECT 11.230 -1.560 11.510 -1.500 ;
        RECT 12.695 -1.555 16.160 -1.500 ;
        RECT 4.980 -1.775 5.300 -1.740 ;
        RECT 5.660 -1.775 5.890 -1.680 ;
        RECT 6.130 -1.770 6.360 -1.680 ;
        RECT 4.980 -1.965 5.890 -1.775 ;
        RECT 4.980 -2.000 5.300 -1.965 ;
        RECT 5.660 -2.100 5.890 -1.965 ;
        RECT 6.120 -1.980 7.360 -1.770 ;
        RECT 6.130 -2.100 6.360 -1.980 ;
        RECT 5.865 -2.315 6.155 -2.260 ;
        RECT 3.750 -2.490 6.155 -2.315 ;
        RECT 3.750 -2.525 6.135 -2.490 ;
        RECT 7.150 -2.745 7.360 -1.980 ;
        RECT 6.345 -2.760 7.360 -2.745 ;
        RECT 5.150 -2.955 7.360 -2.760 ;
        RECT 5.150 -3.480 6.900 -2.955 ;
        RECT 3.140 -7.120 5.740 -6.840 ;
        RECT 6.000 -8.110 6.310 -3.480 ;
        RECT 12.160 -4.180 12.420 -4.145 ;
        RECT 11.305 -4.430 12.420 -4.180 ;
        RECT 11.305 -4.730 11.555 -4.430 ;
        RECT 12.160 -4.465 12.420 -4.430 ;
        RECT 10.540 -4.980 11.560 -4.730 ;
        RECT 12.695 -4.805 12.865 -1.555 ;
        RECT 15.310 -2.160 15.630 -1.900 ;
        RECT 13.210 -4.180 13.530 -4.175 ;
        RECT 13.210 -4.430 14.750 -4.180 ;
        RECT 13.210 -4.435 13.530 -4.430 ;
        RECT 14.445 -4.440 14.735 -4.430 ;
        RECT 14.240 -4.805 14.470 -4.600 ;
        RECT 12.695 -4.975 14.470 -4.805 ;
        RECT 6.810 -6.840 7.085 -6.810 ;
        RECT 6.810 -7.115 10.305 -6.840 ;
        RECT 6.810 -7.145 7.085 -7.115 ;
        RECT 10.540 -8.110 10.790 -4.980 ;
        RECT 11.305 -5.235 11.555 -4.980 ;
        RECT 14.240 -5.020 14.470 -4.975 ;
        RECT 14.710 -4.770 14.940 -4.600 ;
        RECT 15.380 -4.770 15.560 -2.160 ;
        RECT 14.710 -4.950 15.560 -4.770 ;
        RECT 14.710 -5.020 14.940 -4.950 ;
        RECT 15.380 -5.140 15.560 -4.950 ;
        RECT 14.445 -5.235 14.735 -5.180 ;
        RECT 11.305 -5.485 14.765 -5.235 ;
        RECT 15.040 -5.320 15.560 -5.140 ;
        RECT 15.040 -5.690 15.220 -5.320 ;
        RECT 13.810 -5.920 15.370 -5.690 ;
        RECT 20.240 -6.200 20.420 -0.620 ;
        RECT 22.160 -3.470 22.340 0.050 ;
        RECT 37.825 0.215 38.645 0.220 ;
        RECT 25.180 -3.070 26.210 -2.890 ;
        RECT 25.180 -3.470 25.360 -3.070 ;
        RECT 25.905 -3.130 26.195 -3.070 ;
        RECT 25.700 -3.390 25.930 -3.290 ;
        RECT 26.170 -3.390 26.400 -3.290 ;
        RECT 26.740 -3.390 26.970 -2.530 ;
        RECT 22.160 -3.650 25.360 -3.470 ;
        RECT 25.670 -3.580 29.340 -3.390 ;
        RECT 25.040 -3.900 25.220 -3.650 ;
        RECT 25.700 -3.710 25.930 -3.580 ;
        RECT 26.170 -3.710 26.400 -3.580 ;
        RECT 25.905 -3.900 26.195 -3.870 ;
        RECT 25.040 -4.080 26.195 -3.900 ;
        RECT 25.905 -4.100 26.195 -4.080 ;
        RECT 26.740 -4.470 26.970 -3.580 ;
        RECT 29.150 -5.965 29.340 -3.580 ;
        RECT 37.825 -5.965 38.015 0.215 ;
        RECT 29.150 -6.155 38.015 -5.965 ;
        RECT 20.170 -6.460 20.490 -6.200 ;
        RECT 11.090 -6.840 11.365 -6.810 ;
        RECT 11.090 -7.115 21.945 -6.840 ;
        RECT 11.090 -7.145 11.365 -7.115 ;
        RECT 20.170 -7.740 20.490 -7.480 ;
        RECT 1.165 -8.160 20.040 -8.110 ;
        RECT 20.240 -8.160 20.420 -7.740 ;
        RECT 1.165 -8.410 20.550 -8.160 ;
        RECT 1.165 -8.420 12.080 -8.410 ;
        RECT 14.200 -8.420 20.550 -8.410 ;
        RECT -31.175 -10.865 5.705 -10.535 ;
        RECT 5.375 -17.905 5.705 -10.865 ;
        RECT 9.940 -16.330 10.380 -8.420 ;
        RECT 16.715 -10.740 17.025 -8.420 ;
        RECT 17.690 -9.915 17.880 -9.880 ;
        RECT 21.670 -9.915 21.945 -7.115 ;
        RECT 29.150 -9.130 29.340 -6.155 ;
        RECT 29.115 -9.450 29.375 -9.130 ;
        RECT 17.690 -10.105 33.375 -9.915 ;
        RECT 16.715 -11.085 17.390 -10.740 ;
        RECT 16.810 -12.380 17.390 -11.085 ;
        RECT 17.690 -11.375 17.880 -10.105 ;
        RECT 21.670 -10.165 21.945 -10.105 ;
        RECT 29.085 -10.620 29.405 -10.360 ;
        RECT 29.150 -11.170 29.340 -10.620 ;
        RECT 17.670 -11.665 17.900 -11.375 ;
        RECT 26.905 -11.400 32.975 -11.170 ;
        RECT 33.185 -11.375 33.375 -10.105 ;
        RECT 40.950 -10.600 41.390 5.050 ;
        RECT 44.390 3.490 44.790 3.830 ;
        RECT 44.420 -8.135 44.760 3.490 ;
        RECT 51.405 0.310 51.735 8.925 ;
        RECT 84.005 2.945 84.295 18.365 ;
        RECT 85.470 18.020 86.470 18.365 ;
        RECT 85.790 17.290 85.990 18.020 ;
        RECT 87.130 4.260 87.470 25.010 ;
        RECT 91.160 24.830 92.160 25.010 ;
        RECT 91.580 24.440 91.880 24.830 ;
        RECT 91.150 23.090 92.150 24.440 ;
        RECT 90.150 22.905 90.470 22.920 ;
        RECT 90.750 22.905 92.560 23.090 ;
        RECT 90.150 22.675 92.560 22.905 ;
        RECT 90.150 22.660 90.470 22.675 ;
        RECT 90.750 22.220 92.560 22.675 ;
        RECT 91.550 21.910 91.840 21.920 ;
        RECT 89.560 21.650 91.890 21.910 ;
        RECT 88.250 18.720 89.250 19.020 ;
        RECT 87.830 18.550 89.250 18.720 ;
        RECT 89.560 18.760 89.820 21.650 ;
        RECT 90.150 21.360 90.470 21.375 ;
        RECT 91.360 21.360 91.590 21.485 ;
        RECT 90.150 21.130 91.590 21.360 ;
        RECT 90.150 21.115 90.470 21.130 ;
        RECT 91.360 18.985 91.590 21.130 ;
        RECT 91.800 20.230 92.030 21.485 ;
        RECT 91.800 20.020 93.310 20.230 ;
        RECT 91.800 18.985 92.030 20.020 ;
        RECT 91.550 18.760 91.840 18.780 ;
        RECT 89.560 18.550 91.890 18.760 ;
        RECT 87.830 18.500 91.890 18.550 ;
        RECT 87.830 18.480 89.840 18.500 ;
        RECT 88.250 18.260 89.840 18.480 ;
        RECT 88.250 17.990 89.250 18.260 ;
        RECT 89.560 16.740 89.820 18.260 ;
        RECT 93.055 18.130 93.265 20.020 ;
        RECT 93.050 17.840 93.835 18.130 ;
        RECT 94.045 17.875 94.315 29.535 ;
        RECT 106.165 28.850 106.345 29.950 ;
        RECT 108.315 29.820 109.795 30.820 ;
        RECT 109.965 30.400 110.165 31.510 ;
        RECT 124.890 31.495 128.385 31.785 ;
        RECT 109.950 30.140 112.880 30.400 ;
        RECT 108.315 29.680 108.905 29.820 ;
        RECT 109.965 29.090 110.165 30.140 ;
        RECT 108.215 29.080 110.165 29.090 ;
        RECT 102.110 28.670 106.345 28.850 ;
        RECT 108.005 28.890 110.165 29.080 ;
        RECT 108.005 28.740 108.275 28.890 ;
        RECT 96.425 21.880 97.425 22.910 ;
        RECT 96.755 21.260 97.005 21.880 ;
        RECT 98.435 21.260 98.695 21.280 ;
        RECT 95.225 20.960 98.705 21.260 ;
        RECT 95.265 19.520 95.525 20.960 ;
        RECT 97.695 19.860 97.955 20.180 ;
        RECT 97.725 19.710 97.925 19.860 ;
        RECT 95.265 19.230 95.555 19.520 ;
        RECT 95.760 19.480 98.260 19.710 ;
        RECT 95.265 19.170 95.525 19.230 ;
        RECT 95.760 19.040 98.260 19.270 ;
        RECT 98.435 19.190 98.695 20.960 ;
        RECT 99.045 20.710 99.305 20.770 ;
        RECT 99.045 20.510 100.885 20.710 ;
        RECT 99.045 20.450 99.305 20.510 ;
        RECT 98.960 19.910 99.480 20.080 ;
        RECT 96.835 17.885 97.025 19.040 ;
        RECT 98.960 18.890 100.270 19.910 ;
        RECT 98.960 18.510 99.480 18.890 ;
        RECT 94.580 17.875 97.030 17.885 ;
        RECT 90.580 17.625 90.900 17.650 ;
        RECT 93.055 17.625 93.265 17.840 ;
        RECT 90.580 17.415 93.265 17.625 ;
        RECT 94.045 17.620 97.030 17.875 ;
        RECT 100.685 17.850 100.885 20.510 ;
        RECT 102.110 17.850 102.290 28.670 ;
        RECT 104.425 28.000 105.165 28.250 ;
        RECT 103.635 27.000 105.165 28.000 ;
        RECT 106.165 27.780 106.345 28.670 ;
        RECT 104.425 26.660 105.165 27.000 ;
        RECT 105.425 27.590 105.665 27.600 ;
        RECT 105.425 27.300 105.695 27.590 ;
        RECT 105.855 27.550 106.855 27.780 ;
        RECT 105.425 26.200 105.665 27.300 ;
        RECT 105.855 27.110 106.855 27.340 ;
        RECT 106.995 27.140 107.255 27.640 ;
        RECT 106.265 26.920 106.465 27.110 ;
        RECT 108.025 26.920 108.225 28.740 ;
        RECT 106.265 26.720 108.225 26.920 ;
        RECT 106.965 26.200 107.285 26.210 ;
        RECT 105.425 25.960 107.285 26.200 ;
        RECT 105.705 24.630 106.705 25.960 ;
        RECT 106.965 25.950 107.285 25.960 ;
        RECT 104.725 22.900 105.725 23.940 ;
        RECT 110.125 22.900 111.125 24.130 ;
        RECT 103.875 22.635 104.195 22.660 ;
        RECT 104.445 22.635 106.185 22.900 ;
        RECT 109.825 22.700 111.555 22.900 ;
        RECT 103.875 22.425 106.185 22.635 ;
        RECT 109.555 22.440 111.555 22.700 ;
        RECT 103.875 22.400 104.195 22.425 ;
        RECT 104.445 21.960 106.185 22.425 ;
        RECT 109.825 22.040 111.555 22.440 ;
        RECT 105.055 21.700 105.345 21.720 ;
        RECT 103.375 21.460 105.345 21.700 ;
        RECT 108.620 21.480 110.880 21.780 ;
        RECT 103.375 18.590 103.655 21.460 ;
        RECT 103.875 21.100 104.195 21.125 ;
        RECT 104.865 21.100 105.095 21.285 ;
        RECT 103.875 20.890 105.095 21.100 ;
        RECT 103.875 20.865 104.195 20.890 ;
        RECT 104.865 18.785 105.095 20.890 ;
        RECT 105.305 19.900 105.535 21.285 ;
        RECT 105.305 19.740 106.535 19.900 ;
        RECT 105.305 18.785 105.535 19.740 ;
        RECT 103.375 18.350 105.395 18.590 ;
        RECT 103.375 17.850 103.655 18.350 ;
        RECT 106.375 18.030 106.535 19.740 ;
        RECT 108.620 18.600 108.920 21.480 ;
        RECT 110.315 21.010 110.545 21.275 ;
        RECT 109.085 20.990 109.405 21.000 ;
        RECT 109.595 20.990 110.545 21.010 ;
        RECT 109.085 20.770 110.545 20.990 ;
        RECT 109.085 20.750 109.845 20.770 ;
        RECT 109.085 20.740 109.405 20.750 ;
        RECT 110.315 18.775 110.545 20.770 ;
        RECT 110.755 19.780 110.985 21.275 ;
        RECT 110.755 19.570 112.200 19.780 ;
        RECT 110.755 18.775 110.985 19.570 ;
        RECT 108.620 18.300 110.840 18.600 ;
        RECT 108.620 18.120 108.920 18.300 ;
        RECT 108.500 18.090 108.920 18.120 ;
        RECT 107.200 18.030 108.920 18.090 ;
        RECT 94.045 17.605 94.755 17.620 ;
        RECT 90.580 17.390 90.900 17.415 ;
        RECT 95.120 17.110 95.770 17.410 ;
        RECT 89.560 16.480 91.900 16.740 ;
        RECT 89.580 15.150 89.840 16.480 ;
        RECT 91.530 16.470 91.820 16.480 ;
        RECT 90.580 15.895 90.900 15.920 ;
        RECT 91.340 15.895 91.570 16.310 ;
        RECT 90.580 15.685 91.570 15.895 ;
        RECT 90.580 15.660 90.900 15.685 ;
        RECT 91.340 15.310 91.570 15.685 ;
        RECT 91.780 15.900 92.010 16.310 ;
        RECT 94.290 16.110 95.770 17.110 ;
        RECT 96.835 16.850 97.025 17.620 ;
        RECT 100.670 17.610 103.655 17.850 ;
        RECT 106.365 17.840 108.920 18.030 ;
        RECT 106.365 17.790 107.715 17.840 ;
        RECT 98.895 17.410 100.885 17.610 ;
        RECT 102.110 17.600 102.290 17.610 ;
        RECT 91.780 15.680 92.770 15.900 ;
        RECT 91.780 15.310 92.010 15.680 ;
        RECT 89.580 14.890 91.840 15.150 ;
        RECT 92.540 14.640 92.760 15.680 ;
        RECT 95.120 15.640 95.770 16.110 ;
        RECT 96.060 16.660 96.250 16.685 ;
        RECT 96.060 16.370 96.295 16.660 ;
        RECT 96.455 16.620 97.455 16.850 ;
        RECT 96.060 15.215 96.250 16.370 ;
        RECT 96.455 16.180 97.455 16.410 ;
        RECT 97.615 16.390 97.845 16.660 ;
        RECT 96.885 15.810 97.085 16.180 ;
        RECT 97.600 16.070 97.860 16.390 ;
        RECT 98.895 16.150 99.095 17.410 ;
        RECT 103.375 16.970 103.655 17.610 ;
        RECT 104.335 17.640 104.655 17.690 ;
        RECT 106.375 17.640 106.535 17.790 ;
        RECT 104.335 17.480 106.535 17.640 ;
        RECT 107.200 17.610 107.715 17.790 ;
        RECT 104.335 17.430 104.655 17.480 ;
        RECT 103.375 16.730 105.405 16.970 ;
        RECT 103.395 16.690 105.405 16.730 ;
        RECT 98.895 16.060 99.105 16.150 ;
        RECT 98.905 15.810 99.105 16.060 ;
        RECT 96.885 15.610 99.105 15.810 ;
        RECT 103.405 15.370 103.695 16.690 ;
        RECT 105.085 16.680 105.375 16.690 ;
        RECT 104.335 16.180 104.655 16.230 ;
        RECT 104.895 16.180 105.125 16.520 ;
        RECT 104.335 16.020 105.125 16.180 ;
        RECT 104.335 15.970 104.655 16.020 ;
        RECT 104.895 15.520 105.125 16.020 ;
        RECT 105.335 16.130 105.565 16.520 ;
        RECT 105.335 15.930 106.225 16.130 ;
        RECT 105.335 15.520 105.565 15.930 ;
        RECT 97.600 15.215 97.860 15.280 ;
        RECT 96.060 15.025 97.860 15.215 ;
        RECT 103.405 15.090 105.425 15.370 ;
        RECT 90.770 14.320 92.760 14.640 ;
        RECT 96.855 14.400 97.075 15.025 ;
        RECT 97.600 14.960 97.860 15.025 ;
        RECT 105.965 14.840 106.165 15.930 ;
        RECT 104.395 14.640 106.165 14.840 ;
        RECT 90.770 14.060 92.550 14.320 ;
        RECT 104.395 14.180 106.155 14.640 ;
        RECT 91.150 13.070 92.150 14.060 ;
        RECT 104.725 13.440 105.725 14.180 ;
        RECT 91.510 12.740 91.790 13.070 ;
        RECT 88.450 12.230 88.890 12.260 ;
        RECT 91.130 12.230 92.130 12.740 ;
        RECT 107.465 12.515 107.715 17.610 ;
        RECT 108.620 16.590 108.920 17.840 ;
        RECT 111.985 17.880 112.195 19.570 ;
        RECT 112.620 17.880 112.880 30.140 ;
        RECT 124.890 29.710 125.180 31.495 ;
        RECT 127.315 30.740 130.915 30.960 ;
        RECT 127.315 29.900 127.535 30.740 ;
        RECT 128.715 30.110 129.515 30.530 ;
        RECT 124.890 29.420 125.215 29.710 ;
        RECT 125.420 29.670 127.920 29.900 ;
        RECT 124.890 29.375 125.180 29.420 ;
        RECT 125.420 29.230 127.920 29.460 ;
        RECT 128.065 29.390 128.355 30.070 ;
        RECT 126.455 28.260 126.655 29.230 ;
        RECT 128.715 29.110 130.375 30.110 ;
        RECT 130.695 29.915 130.915 30.740 ;
        RECT 130.695 29.645 132.465 29.915 ;
        RECT 128.715 28.830 129.515 29.110 ;
        RECT 121.300 28.060 126.655 28.260 ;
        RECT 130.695 28.210 130.915 29.645 ;
        RECT 116.415 21.840 116.725 22.480 ;
        RECT 115.015 21.540 118.465 21.840 ;
        RECT 115.015 19.680 115.315 21.540 ;
        RECT 117.715 21.030 120.485 21.210 ;
        RECT 117.715 20.190 117.895 21.030 ;
        RECT 118.705 20.440 119.565 20.720 ;
        RECT 115.460 19.960 117.960 20.190 ;
        RECT 115.460 19.520 117.960 19.750 ;
        RECT 118.135 19.710 118.435 20.270 ;
        RECT 116.365 18.425 116.545 19.520 ;
        RECT 118.705 19.440 120.145 20.440 ;
        RECT 118.705 19.010 119.565 19.440 ;
        RECT 120.305 18.840 120.485 21.030 ;
        RECT 121.300 18.840 121.500 28.060 ;
        RECT 125.025 27.240 125.435 27.580 ;
        RECT 124.095 26.240 125.435 27.240 ;
        RECT 126.455 27.030 126.655 28.060 ;
        RECT 128.305 27.990 130.915 28.210 ;
        RECT 125.675 26.840 125.880 26.890 ;
        RECT 125.655 26.550 125.885 26.840 ;
        RECT 126.045 26.800 127.045 27.030 ;
        RECT 125.025 25.820 125.435 26.240 ;
        RECT 125.675 25.530 125.880 26.550 ;
        RECT 126.045 26.360 127.045 26.590 ;
        RECT 126.495 26.080 126.715 26.360 ;
        RECT 127.195 26.250 127.475 26.860 ;
        RECT 128.305 26.080 128.525 27.990 ;
        RECT 126.495 25.860 128.525 26.080 ;
        RECT 125.635 25.250 127.505 25.530 ;
        RECT 126.315 24.610 126.665 25.250 ;
        RECT 122.460 23.010 122.780 23.045 ;
        RECT 123.425 23.040 124.425 24.600 ;
        RECT 123.065 23.010 124.885 23.040 ;
        RECT 122.460 22.820 124.885 23.010 ;
        RECT 128.495 22.990 129.495 24.380 ;
        RECT 128.135 22.980 129.975 22.990 ;
        RECT 122.460 22.785 122.780 22.820 ;
        RECT 123.065 22.350 124.885 22.820 ;
        RECT 127.335 22.720 129.975 22.980 ;
        RECT 128.135 22.130 129.975 22.720 ;
        RECT 122.080 21.800 124.160 22.080 ;
        RECT 122.080 21.130 122.360 21.800 ;
        RECT 126.715 21.690 129.235 21.990 ;
        RECT 122.080 20.500 122.320 21.130 ;
        RECT 122.490 20.895 122.750 20.960 ;
        RECT 123.675 20.895 123.905 21.645 ;
        RECT 122.490 20.705 123.905 20.895 ;
        RECT 122.490 20.640 122.750 20.705 ;
        RECT 122.080 18.920 122.360 20.500 ;
        RECT 123.675 19.145 123.905 20.705 ;
        RECT 124.115 20.440 124.345 21.645 ;
        RECT 126.715 20.550 127.015 21.690 ;
        RECT 128.885 21.620 129.175 21.690 ;
        RECT 128.695 21.030 128.925 21.415 ;
        RECT 127.335 20.770 128.925 21.030 ;
        RECT 124.115 20.190 125.425 20.440 ;
        RECT 126.715 20.250 127.745 20.550 ;
        RECT 124.115 19.145 124.345 20.190 ;
        RECT 123.865 18.920 124.155 18.940 ;
        RECT 122.080 18.840 124.230 18.920 ;
        RECT 120.295 18.660 124.230 18.840 ;
        RECT 118.525 18.640 124.230 18.660 ;
        RECT 118.525 18.610 122.430 18.640 ;
        RECT 118.525 18.480 120.485 18.610 ;
        RECT 111.985 17.620 112.880 17.880 ;
        RECT 113.725 18.175 116.575 18.425 ;
        RECT 109.800 17.495 110.120 17.520 ;
        RECT 111.985 17.495 112.195 17.620 ;
        RECT 109.800 17.285 112.195 17.495 ;
        RECT 109.800 17.260 110.120 17.285 ;
        RECT 108.620 16.290 110.940 16.590 ;
        RECT 108.620 14.980 108.920 16.290 ;
        RECT 109.800 15.815 110.120 15.840 ;
        RECT 110.375 15.815 110.605 16.140 ;
        RECT 109.800 15.605 110.605 15.815 ;
        RECT 109.800 15.580 110.120 15.605 ;
        RECT 110.375 15.140 110.605 15.605 ;
        RECT 110.815 15.770 111.045 16.140 ;
        RECT 110.815 15.530 111.725 15.770 ;
        RECT 110.815 15.140 111.045 15.530 ;
        RECT 108.620 14.680 110.930 14.980 ;
        RECT 111.485 14.440 111.725 15.530 ;
        RECT 109.750 14.110 111.725 14.440 ;
        RECT 109.750 13.840 111.640 14.110 ;
        RECT 110.360 13.020 111.360 13.840 ;
        RECT 113.725 12.515 113.975 18.175 ;
        RECT 114.995 17.550 115.585 18.000 ;
        RECT 114.255 16.550 115.585 17.550 ;
        RECT 116.365 17.430 116.545 18.175 ;
        RECT 114.995 16.200 115.585 16.550 ;
        RECT 115.845 15.910 116.095 17.270 ;
        RECT 116.255 17.200 117.255 17.430 ;
        RECT 117.425 17.240 117.665 17.250 ;
        RECT 116.255 16.760 117.255 16.990 ;
        RECT 117.415 16.950 117.665 17.240 ;
        RECT 116.645 16.360 116.825 16.760 ;
        RECT 117.415 16.630 117.675 16.950 ;
        RECT 117.425 16.600 117.665 16.630 ;
        RECT 118.525 16.360 118.705 18.480 ;
        RECT 116.645 16.180 118.705 16.360 ;
        RECT 122.080 17.260 122.360 18.610 ;
        RECT 125.170 18.560 125.420 20.190 ;
        RECT 127.445 18.740 127.745 20.250 ;
        RECT 128.695 18.915 128.925 20.770 ;
        RECT 129.135 20.150 129.365 21.415 ;
        RECT 129.135 19.890 130.635 20.150 ;
        RECT 129.135 18.915 129.365 19.890 ;
        RECT 127.435 18.630 129.255 18.740 ;
        RECT 126.695 18.560 129.255 18.630 ;
        RECT 125.170 18.440 129.255 18.560 ;
        RECT 125.170 18.360 127.745 18.440 ;
        RECT 125.170 18.330 126.945 18.360 ;
        RECT 122.865 18.075 123.185 18.080 ;
        RECT 125.170 18.075 125.420 18.330 ;
        RECT 122.865 17.825 125.420 18.075 ;
        RECT 122.865 17.820 123.185 17.825 ;
        RECT 122.080 16.980 124.210 17.260 ;
        RECT 115.835 15.650 116.095 15.910 ;
        RECT 117.385 15.720 117.705 15.980 ;
        RECT 115.835 15.500 116.075 15.650 ;
        RECT 117.425 15.500 117.665 15.720 ;
        RECT 115.835 15.260 117.665 15.500 ;
        RECT 122.080 15.600 122.360 16.980 ;
        RECT 123.895 16.940 124.185 16.980 ;
        RECT 122.895 16.385 123.155 16.420 ;
        RECT 123.705 16.385 123.935 16.780 ;
        RECT 122.895 16.135 123.935 16.385 ;
        RECT 124.145 16.350 124.375 16.780 ;
        RECT 122.895 16.100 123.155 16.135 ;
        RECT 123.705 15.780 123.935 16.135 ;
        RECT 124.105 16.070 125.215 16.350 ;
        RECT 124.145 15.780 124.375 16.070 ;
        RECT 123.895 15.600 124.185 15.620 ;
        RECT 122.080 15.390 124.185 15.600 ;
        RECT 122.080 15.320 124.170 15.390 ;
        RECT 115.965 14.920 117.515 15.260 ;
        RECT 124.935 15.130 125.215 16.070 ;
        RECT 116.275 14.040 117.275 14.920 ;
        RECT 123.095 14.670 125.215 15.130 ;
        RECT 123.095 14.350 124.935 14.670 ;
        RECT 123.775 13.550 124.775 14.350 ;
        RECT 107.465 12.265 113.975 12.515 ;
        RECT 126.180 12.690 126.400 18.330 ;
        RECT 127.435 16.940 127.735 18.360 ;
        RECT 130.375 18.320 130.635 19.890 ;
        RECT 132.195 18.320 132.465 29.645 ;
        RECT 132.895 18.320 133.165 36.265 ;
        RECT 140.465 32.935 140.735 38.120 ;
        RECT 152.030 36.165 155.530 36.235 ;
        RECT 152.030 35.965 182.100 36.165 ;
        RECT 140.465 32.605 141.815 32.935 ;
        RECT 140.465 24.070 140.735 32.605 ;
        RECT 152.030 29.435 152.300 35.965 ;
        RECT 155.155 35.895 182.100 35.965 ;
        RECT 155.020 31.890 155.330 32.320 ;
        RECT 156.695 31.890 156.955 31.950 ;
        RECT 153.570 31.690 156.955 31.890 ;
        RECT 175.120 31.840 176.120 32.870 ;
        RECT 153.570 30.060 153.770 31.690 ;
        RECT 155.020 31.680 155.330 31.690 ;
        RECT 156.695 31.630 156.955 31.690 ;
        RECT 175.410 31.415 175.730 31.840 ;
        RECT 155.780 31.140 159.100 31.340 ;
        RECT 155.780 30.250 155.980 31.140 ;
        RECT 157.250 30.450 157.840 30.760 ;
        RECT 153.570 29.770 153.800 30.060 ;
        RECT 154.005 30.020 156.505 30.250 ;
        RECT 156.695 30.150 156.955 30.450 ;
        RECT 153.570 29.760 153.770 29.770 ;
        RECT 154.005 29.580 156.505 29.810 ;
        RECT 156.660 29.720 156.990 30.150 ;
        RECT 142.980 29.165 152.300 29.435 ;
        RECT 140.085 22.720 141.085 24.070 ;
        RECT 139.085 22.535 139.405 22.550 ;
        RECT 139.685 22.535 141.495 22.720 ;
        RECT 139.085 22.305 141.495 22.535 ;
        RECT 139.085 22.290 139.405 22.305 ;
        RECT 139.685 21.850 141.495 22.305 ;
        RECT 140.485 21.540 140.775 21.550 ;
        RECT 138.495 21.280 140.825 21.540 ;
        RECT 130.375 18.050 134.835 18.320 ;
        RECT 137.185 18.180 138.185 18.650 ;
        RECT 138.495 18.390 138.755 21.280 ;
        RECT 139.085 20.990 139.405 21.005 ;
        RECT 140.295 20.990 140.525 21.115 ;
        RECT 139.085 20.760 140.525 20.990 ;
        RECT 139.085 20.745 139.405 20.760 ;
        RECT 140.295 18.615 140.525 20.760 ;
        RECT 140.735 19.860 140.965 21.115 ;
        RECT 140.735 19.650 142.245 19.860 ;
        RECT 140.735 18.615 140.965 19.650 ;
        RECT 140.485 18.390 140.775 18.410 ;
        RECT 138.495 18.180 140.825 18.390 ;
        RECT 137.185 18.140 140.825 18.180 ;
        RECT 137.010 18.130 140.825 18.140 ;
        RECT 130.375 17.840 130.635 18.050 ;
        RECT 128.005 17.580 130.635 17.840 ;
        RECT 137.010 17.890 138.775 18.130 ;
        RECT 137.010 17.620 138.185 17.890 ;
        RECT 137.010 17.180 137.230 17.620 ;
        RECT 131.610 16.960 137.230 17.180 ;
        RECT 127.365 16.870 129.195 16.940 ;
        RECT 127.365 16.640 129.205 16.870 ;
        RECT 127.435 15.320 127.735 16.640 ;
        RECT 128.725 16.100 128.955 16.480 ;
        RECT 128.005 15.840 128.955 16.100 ;
        RECT 128.725 15.480 128.955 15.840 ;
        RECT 129.165 15.750 129.395 16.480 ;
        RECT 129.165 15.560 130.065 15.750 ;
        RECT 129.165 15.480 129.395 15.560 ;
        RECT 127.435 15.310 128.515 15.320 ;
        RECT 128.915 15.310 129.205 15.320 ;
        RECT 127.435 15.070 129.265 15.310 ;
        RECT 129.875 14.760 130.065 15.560 ;
        RECT 128.105 14.465 130.065 14.760 ;
        RECT 128.105 14.130 130.005 14.465 ;
        RECT 128.605 12.950 129.605 14.130 ;
        RECT 131.610 12.690 131.830 16.960 ;
        RECT 138.495 16.370 138.755 17.890 ;
        RECT 141.990 17.760 142.200 19.650 ;
        RECT 141.985 17.470 142.770 17.760 ;
        RECT 142.980 17.505 143.250 29.165 ;
        RECT 155.100 28.480 155.280 29.580 ;
        RECT 157.250 29.450 158.730 30.450 ;
        RECT 158.900 30.030 159.100 31.140 ;
        RECT 173.825 31.125 177.320 31.415 ;
        RECT 158.885 29.770 161.815 30.030 ;
        RECT 157.250 29.310 157.840 29.450 ;
        RECT 158.900 28.720 159.100 29.770 ;
        RECT 157.150 28.710 159.100 28.720 ;
        RECT 151.045 28.300 155.280 28.480 ;
        RECT 156.940 28.520 159.100 28.710 ;
        RECT 156.940 28.370 157.210 28.520 ;
        RECT 145.360 21.510 146.360 22.540 ;
        RECT 145.690 20.890 145.940 21.510 ;
        RECT 147.370 20.890 147.630 20.910 ;
        RECT 144.160 20.590 147.640 20.890 ;
        RECT 144.200 19.150 144.460 20.590 ;
        RECT 146.630 19.490 146.890 19.810 ;
        RECT 146.660 19.340 146.860 19.490 ;
        RECT 144.200 18.860 144.490 19.150 ;
        RECT 144.695 19.110 147.195 19.340 ;
        RECT 144.200 18.800 144.460 18.860 ;
        RECT 144.695 18.670 147.195 18.900 ;
        RECT 147.370 18.820 147.630 20.590 ;
        RECT 147.980 20.340 148.240 20.400 ;
        RECT 147.980 20.140 149.820 20.340 ;
        RECT 147.980 20.080 148.240 20.140 ;
        RECT 147.895 19.540 148.415 19.710 ;
        RECT 145.770 17.515 145.960 18.670 ;
        RECT 147.895 18.520 149.205 19.540 ;
        RECT 147.895 18.140 148.415 18.520 ;
        RECT 143.515 17.505 145.965 17.515 ;
        RECT 139.515 17.255 139.835 17.280 ;
        RECT 141.990 17.255 142.200 17.470 ;
        RECT 139.515 17.045 142.200 17.255 ;
        RECT 142.980 17.250 145.965 17.505 ;
        RECT 149.620 17.480 149.820 20.140 ;
        RECT 151.045 17.480 151.225 28.300 ;
        RECT 153.360 27.630 154.100 27.880 ;
        RECT 152.570 26.630 154.100 27.630 ;
        RECT 155.100 27.410 155.280 28.300 ;
        RECT 153.360 26.290 154.100 26.630 ;
        RECT 154.360 27.220 154.600 27.230 ;
        RECT 154.360 26.930 154.630 27.220 ;
        RECT 154.790 27.180 155.790 27.410 ;
        RECT 154.360 25.830 154.600 26.930 ;
        RECT 154.790 26.740 155.790 26.970 ;
        RECT 155.930 26.770 156.190 27.270 ;
        RECT 155.200 26.550 155.400 26.740 ;
        RECT 156.960 26.550 157.160 28.370 ;
        RECT 155.200 26.350 157.160 26.550 ;
        RECT 155.900 25.830 156.220 25.840 ;
        RECT 154.360 25.590 156.220 25.830 ;
        RECT 154.640 24.260 155.640 25.590 ;
        RECT 155.900 25.580 156.220 25.590 ;
        RECT 153.660 22.530 154.660 23.570 ;
        RECT 159.060 22.530 160.060 23.760 ;
        RECT 152.810 22.265 153.130 22.290 ;
        RECT 153.380 22.265 155.120 22.530 ;
        RECT 158.760 22.330 160.490 22.530 ;
        RECT 152.810 22.055 155.120 22.265 ;
        RECT 158.490 22.070 160.490 22.330 ;
        RECT 152.810 22.030 153.130 22.055 ;
        RECT 153.380 21.590 155.120 22.055 ;
        RECT 158.760 21.670 160.490 22.070 ;
        RECT 153.990 21.330 154.280 21.350 ;
        RECT 152.310 21.090 154.280 21.330 ;
        RECT 157.555 21.110 159.815 21.410 ;
        RECT 152.310 18.220 152.590 21.090 ;
        RECT 152.810 20.730 153.130 20.755 ;
        RECT 153.800 20.730 154.030 20.915 ;
        RECT 152.810 20.520 154.030 20.730 ;
        RECT 152.810 20.495 153.130 20.520 ;
        RECT 153.800 18.415 154.030 20.520 ;
        RECT 154.240 19.530 154.470 20.915 ;
        RECT 154.240 19.370 155.470 19.530 ;
        RECT 154.240 18.415 154.470 19.370 ;
        RECT 152.310 17.980 154.330 18.220 ;
        RECT 152.310 17.480 152.590 17.980 ;
        RECT 155.310 17.660 155.470 19.370 ;
        RECT 157.555 18.230 157.855 21.110 ;
        RECT 159.250 20.640 159.480 20.905 ;
        RECT 158.020 20.620 158.340 20.630 ;
        RECT 158.530 20.620 159.480 20.640 ;
        RECT 158.020 20.400 159.480 20.620 ;
        RECT 158.020 20.380 158.780 20.400 ;
        RECT 158.020 20.370 158.340 20.380 ;
        RECT 159.250 18.405 159.480 20.400 ;
        RECT 159.690 19.410 159.920 20.905 ;
        RECT 159.690 19.200 161.135 19.410 ;
        RECT 159.690 18.405 159.920 19.200 ;
        RECT 157.555 17.930 159.775 18.230 ;
        RECT 157.555 17.750 157.855 17.930 ;
        RECT 157.435 17.720 157.855 17.750 ;
        RECT 156.135 17.660 157.855 17.720 ;
        RECT 142.980 17.235 143.690 17.250 ;
        RECT 139.515 17.020 139.835 17.045 ;
        RECT 144.055 16.740 144.705 17.040 ;
        RECT 138.495 16.110 140.835 16.370 ;
        RECT 138.515 14.780 138.775 16.110 ;
        RECT 140.465 16.100 140.755 16.110 ;
        RECT 139.515 15.525 139.835 15.550 ;
        RECT 140.275 15.525 140.505 15.940 ;
        RECT 139.515 15.315 140.505 15.525 ;
        RECT 139.515 15.290 139.835 15.315 ;
        RECT 140.275 14.940 140.505 15.315 ;
        RECT 140.715 15.530 140.945 15.940 ;
        RECT 143.225 15.740 144.705 16.740 ;
        RECT 145.770 16.480 145.960 17.250 ;
        RECT 149.605 17.240 152.590 17.480 ;
        RECT 155.300 17.470 157.855 17.660 ;
        RECT 155.300 17.420 156.650 17.470 ;
        RECT 147.830 17.040 149.820 17.240 ;
        RECT 151.045 17.230 151.225 17.240 ;
        RECT 140.715 15.310 141.705 15.530 ;
        RECT 140.715 14.940 140.945 15.310 ;
        RECT 138.515 14.520 140.775 14.780 ;
        RECT 141.475 14.270 141.695 15.310 ;
        RECT 144.055 15.270 144.705 15.740 ;
        RECT 144.995 16.290 145.185 16.315 ;
        RECT 144.995 16.000 145.230 16.290 ;
        RECT 145.390 16.250 146.390 16.480 ;
        RECT 144.995 14.845 145.185 16.000 ;
        RECT 145.390 15.810 146.390 16.040 ;
        RECT 146.550 16.020 146.780 16.290 ;
        RECT 145.820 15.440 146.020 15.810 ;
        RECT 146.535 15.700 146.795 16.020 ;
        RECT 147.830 15.780 148.030 17.040 ;
        RECT 152.310 16.600 152.590 17.240 ;
        RECT 153.270 17.270 153.590 17.320 ;
        RECT 155.310 17.270 155.470 17.420 ;
        RECT 153.270 17.110 155.470 17.270 ;
        RECT 156.135 17.240 156.650 17.420 ;
        RECT 153.270 17.060 153.590 17.110 ;
        RECT 152.310 16.360 154.340 16.600 ;
        RECT 152.330 16.320 154.340 16.360 ;
        RECT 147.830 15.690 148.040 15.780 ;
        RECT 147.840 15.440 148.040 15.690 ;
        RECT 145.820 15.240 148.040 15.440 ;
        RECT 152.340 15.000 152.630 16.320 ;
        RECT 154.020 16.310 154.310 16.320 ;
        RECT 153.270 15.810 153.590 15.860 ;
        RECT 153.830 15.810 154.060 16.150 ;
        RECT 153.270 15.650 154.060 15.810 ;
        RECT 153.270 15.600 153.590 15.650 ;
        RECT 153.830 15.150 154.060 15.650 ;
        RECT 154.270 15.760 154.500 16.150 ;
        RECT 154.270 15.560 155.160 15.760 ;
        RECT 154.270 15.150 154.500 15.560 ;
        RECT 146.535 14.845 146.795 14.910 ;
        RECT 144.995 14.655 146.795 14.845 ;
        RECT 152.340 14.720 154.360 15.000 ;
        RECT 139.705 13.950 141.695 14.270 ;
        RECT 145.790 14.030 146.010 14.655 ;
        RECT 146.535 14.590 146.795 14.655 ;
        RECT 154.900 14.470 155.100 15.560 ;
        RECT 153.330 14.270 155.100 14.470 ;
        RECT 139.705 13.690 141.485 13.950 ;
        RECT 153.330 13.810 155.090 14.270 ;
        RECT 140.085 12.700 141.085 13.690 ;
        RECT 153.660 13.070 154.660 13.810 ;
        RECT 126.180 12.470 131.830 12.690 ;
        RECT 88.450 11.790 92.130 12.230 ;
        RECT 88.450 11.760 88.890 11.790 ;
        RECT 91.130 11.740 92.130 11.790 ;
        RECT 91.460 10.940 91.780 11.740 ;
        RECT 140.490 10.940 140.810 12.700 ;
        RECT 156.400 12.145 156.650 17.240 ;
        RECT 157.555 16.220 157.855 17.470 ;
        RECT 160.920 17.510 161.130 19.200 ;
        RECT 161.555 17.510 161.815 29.770 ;
        RECT 173.825 29.340 174.115 31.125 ;
        RECT 176.250 30.370 179.850 30.590 ;
        RECT 176.250 29.530 176.470 30.370 ;
        RECT 177.650 29.740 178.450 30.160 ;
        RECT 173.825 29.050 174.150 29.340 ;
        RECT 174.355 29.300 176.855 29.530 ;
        RECT 173.825 29.005 174.115 29.050 ;
        RECT 174.355 28.860 176.855 29.090 ;
        RECT 177.000 29.020 177.290 29.700 ;
        RECT 175.390 27.890 175.590 28.860 ;
        RECT 177.650 28.740 179.310 29.740 ;
        RECT 179.630 29.545 179.850 30.370 ;
        RECT 179.630 29.275 181.400 29.545 ;
        RECT 177.650 28.460 178.450 28.740 ;
        RECT 170.235 27.690 175.590 27.890 ;
        RECT 179.630 27.840 179.850 29.275 ;
        RECT 165.350 21.470 165.660 22.110 ;
        RECT 163.950 21.170 167.400 21.470 ;
        RECT 163.950 19.310 164.250 21.170 ;
        RECT 166.650 20.660 169.420 20.840 ;
        RECT 166.650 19.820 166.830 20.660 ;
        RECT 167.640 20.070 168.500 20.350 ;
        RECT 164.395 19.590 166.895 19.820 ;
        RECT 164.395 19.150 166.895 19.380 ;
        RECT 167.070 19.340 167.370 19.900 ;
        RECT 165.300 18.055 165.480 19.150 ;
        RECT 167.640 19.070 169.080 20.070 ;
        RECT 167.640 18.640 168.500 19.070 ;
        RECT 169.240 18.470 169.420 20.660 ;
        RECT 170.235 18.470 170.435 27.690 ;
        RECT 173.960 26.870 174.370 27.210 ;
        RECT 173.030 25.870 174.370 26.870 ;
        RECT 175.390 26.660 175.590 27.690 ;
        RECT 177.240 27.620 179.850 27.840 ;
        RECT 174.610 26.470 174.815 26.520 ;
        RECT 174.590 26.180 174.820 26.470 ;
        RECT 174.980 26.430 175.980 26.660 ;
        RECT 173.960 25.450 174.370 25.870 ;
        RECT 174.610 25.160 174.815 26.180 ;
        RECT 174.980 25.990 175.980 26.220 ;
        RECT 175.430 25.710 175.650 25.990 ;
        RECT 176.130 25.880 176.410 26.490 ;
        RECT 177.240 25.710 177.460 27.620 ;
        RECT 175.430 25.490 177.460 25.710 ;
        RECT 174.570 24.880 176.440 25.160 ;
        RECT 175.250 24.240 175.600 24.880 ;
        RECT 171.395 22.640 171.715 22.675 ;
        RECT 172.360 22.670 173.360 24.230 ;
        RECT 172.000 22.640 173.820 22.670 ;
        RECT 171.395 22.450 173.820 22.640 ;
        RECT 177.430 22.620 178.430 24.010 ;
        RECT 177.070 22.610 178.910 22.620 ;
        RECT 171.395 22.415 171.715 22.450 ;
        RECT 172.000 21.980 173.820 22.450 ;
        RECT 176.270 22.350 178.910 22.610 ;
        RECT 177.070 21.760 178.910 22.350 ;
        RECT 171.015 21.430 173.095 21.710 ;
        RECT 171.015 20.760 171.295 21.430 ;
        RECT 175.650 21.320 178.170 21.620 ;
        RECT 171.015 20.130 171.255 20.760 ;
        RECT 171.425 20.525 171.685 20.590 ;
        RECT 172.610 20.525 172.840 21.275 ;
        RECT 171.425 20.335 172.840 20.525 ;
        RECT 171.425 20.270 171.685 20.335 ;
        RECT 171.015 18.550 171.295 20.130 ;
        RECT 172.610 18.775 172.840 20.335 ;
        RECT 173.050 20.070 173.280 21.275 ;
        RECT 175.650 20.180 175.950 21.320 ;
        RECT 177.820 21.250 178.110 21.320 ;
        RECT 177.630 20.660 177.860 21.045 ;
        RECT 176.270 20.400 177.860 20.660 ;
        RECT 173.050 19.820 174.360 20.070 ;
        RECT 175.650 19.880 176.680 20.180 ;
        RECT 173.050 18.775 173.280 19.820 ;
        RECT 172.800 18.550 173.090 18.570 ;
        RECT 171.015 18.470 173.165 18.550 ;
        RECT 169.230 18.290 173.165 18.470 ;
        RECT 167.460 18.270 173.165 18.290 ;
        RECT 167.460 18.240 171.365 18.270 ;
        RECT 167.460 18.110 169.420 18.240 ;
        RECT 160.920 17.250 161.815 17.510 ;
        RECT 162.660 17.805 165.510 18.055 ;
        RECT 158.735 17.125 159.055 17.150 ;
        RECT 160.920 17.125 161.130 17.250 ;
        RECT 158.735 16.915 161.130 17.125 ;
        RECT 158.735 16.890 159.055 16.915 ;
        RECT 157.555 15.920 159.875 16.220 ;
        RECT 157.555 14.610 157.855 15.920 ;
        RECT 158.735 15.445 159.055 15.470 ;
        RECT 159.310 15.445 159.540 15.770 ;
        RECT 158.735 15.235 159.540 15.445 ;
        RECT 158.735 15.210 159.055 15.235 ;
        RECT 159.310 14.770 159.540 15.235 ;
        RECT 159.750 15.400 159.980 15.770 ;
        RECT 159.750 15.160 160.660 15.400 ;
        RECT 159.750 14.770 159.980 15.160 ;
        RECT 157.555 14.310 159.865 14.610 ;
        RECT 160.420 14.070 160.660 15.160 ;
        RECT 158.685 13.740 160.660 14.070 ;
        RECT 158.685 13.470 160.575 13.740 ;
        RECT 159.295 12.650 160.295 13.470 ;
        RECT 162.660 12.145 162.910 17.805 ;
        RECT 163.930 17.180 164.520 17.630 ;
        RECT 163.190 16.180 164.520 17.180 ;
        RECT 165.300 17.060 165.480 17.805 ;
        RECT 163.930 15.830 164.520 16.180 ;
        RECT 164.780 15.540 165.030 16.900 ;
        RECT 165.190 16.830 166.190 17.060 ;
        RECT 166.360 16.870 166.600 16.880 ;
        RECT 165.190 16.390 166.190 16.620 ;
        RECT 166.350 16.580 166.600 16.870 ;
        RECT 165.580 15.990 165.760 16.390 ;
        RECT 166.350 16.260 166.610 16.580 ;
        RECT 166.360 16.230 166.600 16.260 ;
        RECT 167.460 15.990 167.640 18.110 ;
        RECT 165.580 15.810 167.640 15.990 ;
        RECT 171.015 16.890 171.295 18.240 ;
        RECT 174.105 18.190 174.355 19.820 ;
        RECT 176.380 18.370 176.680 19.880 ;
        RECT 177.630 18.545 177.860 20.400 ;
        RECT 178.070 19.780 178.300 21.045 ;
        RECT 178.070 19.520 179.570 19.780 ;
        RECT 178.070 18.545 178.300 19.520 ;
        RECT 176.370 18.260 178.190 18.370 ;
        RECT 175.630 18.190 178.190 18.260 ;
        RECT 174.105 18.070 178.190 18.190 ;
        RECT 174.105 17.990 176.680 18.070 ;
        RECT 174.105 17.960 175.880 17.990 ;
        RECT 171.800 17.705 172.120 17.710 ;
        RECT 174.105 17.705 174.355 17.960 ;
        RECT 171.800 17.455 174.355 17.705 ;
        RECT 171.800 17.450 172.120 17.455 ;
        RECT 171.015 16.610 173.145 16.890 ;
        RECT 164.770 15.280 165.030 15.540 ;
        RECT 166.320 15.350 166.640 15.610 ;
        RECT 164.770 15.130 165.010 15.280 ;
        RECT 166.360 15.130 166.600 15.350 ;
        RECT 164.770 14.890 166.600 15.130 ;
        RECT 171.015 15.230 171.295 16.610 ;
        RECT 172.830 16.570 173.120 16.610 ;
        RECT 171.830 16.015 172.090 16.050 ;
        RECT 172.640 16.015 172.870 16.410 ;
        RECT 171.830 15.765 172.870 16.015 ;
        RECT 173.080 15.980 173.310 16.410 ;
        RECT 171.830 15.730 172.090 15.765 ;
        RECT 172.640 15.410 172.870 15.765 ;
        RECT 173.040 15.700 174.150 15.980 ;
        RECT 173.080 15.410 173.310 15.700 ;
        RECT 172.830 15.230 173.120 15.250 ;
        RECT 171.015 15.020 173.120 15.230 ;
        RECT 171.015 14.950 173.105 15.020 ;
        RECT 164.900 14.550 166.450 14.890 ;
        RECT 173.870 14.760 174.150 15.700 ;
        RECT 165.210 13.670 166.210 14.550 ;
        RECT 172.030 14.300 174.150 14.760 ;
        RECT 172.030 13.980 173.870 14.300 ;
        RECT 172.710 13.180 173.710 13.980 ;
        RECT 156.400 11.895 162.910 12.145 ;
        RECT 175.115 12.320 175.335 17.960 ;
        RECT 176.370 16.570 176.670 17.990 ;
        RECT 179.310 17.950 179.570 19.520 ;
        RECT 181.130 17.950 181.400 29.275 ;
        RECT 181.830 17.950 182.100 35.895 ;
        RECT 179.310 17.680 183.770 17.950 ;
        RECT 179.310 17.470 179.570 17.680 ;
        RECT 176.940 17.210 179.570 17.470 ;
        RECT 180.545 16.590 183.680 16.810 ;
        RECT 176.300 16.500 178.130 16.570 ;
        RECT 176.300 16.270 178.140 16.500 ;
        RECT 176.370 14.950 176.670 16.270 ;
        RECT 177.660 15.730 177.890 16.110 ;
        RECT 176.940 15.470 177.890 15.730 ;
        RECT 177.660 15.110 177.890 15.470 ;
        RECT 178.100 15.380 178.330 16.110 ;
        RECT 178.100 15.190 179.000 15.380 ;
        RECT 178.100 15.110 178.330 15.190 ;
        RECT 176.370 14.940 177.450 14.950 ;
        RECT 177.850 14.940 178.140 14.950 ;
        RECT 176.370 14.700 178.200 14.940 ;
        RECT 178.810 14.390 179.000 15.190 ;
        RECT 177.040 14.095 179.000 14.390 ;
        RECT 177.040 13.760 178.940 14.095 ;
        RECT 177.540 12.580 178.540 13.760 ;
        RECT 180.545 12.320 180.765 16.590 ;
        RECT 183.460 15.750 183.680 16.590 ;
        RECT 175.115 12.100 180.765 12.320 ;
        RECT 91.460 10.620 158.490 10.940 ;
        RECT 118.050 8.615 123.700 8.835 ;
        RECT 115.330 4.440 116.330 4.860 ;
        RECT 114.380 4.345 116.330 4.440 ;
        RECT 118.050 4.345 118.270 8.615 ;
        RECT 120.275 7.175 121.275 8.355 ;
        RECT 119.875 6.840 121.775 7.175 ;
        RECT 119.815 6.545 121.775 6.840 ;
        RECT 119.815 5.745 120.005 6.545 ;
        RECT 120.615 5.995 122.445 6.235 ;
        RECT 120.675 5.985 120.965 5.995 ;
        RECT 121.365 5.985 122.445 5.995 ;
        RECT 120.485 5.745 120.715 5.825 ;
        RECT 119.815 5.555 120.715 5.745 ;
        RECT 120.485 4.825 120.715 5.555 ;
        RECT 120.925 5.465 121.155 5.825 ;
        RECT 120.925 5.205 121.875 5.465 ;
        RECT 120.925 4.825 121.155 5.205 ;
        RECT 122.145 4.665 122.445 5.985 ;
        RECT 120.675 4.435 122.515 4.665 ;
        RECT 120.685 4.365 122.515 4.435 ;
        RECT 87.130 3.920 107.470 4.260 ;
        RECT 84.005 2.655 102.975 2.945 ;
        RECT 55.170 1.825 55.440 1.835 ;
        RECT 62.770 1.825 63.040 1.875 ;
        RECT 70.420 1.825 70.690 1.835 ;
        RECT 78.260 1.825 78.530 1.875 ;
        RECT 86.180 1.825 86.450 1.835 ;
        RECT 93.850 1.825 94.120 1.845 ;
        RECT 53.960 1.555 101.420 1.825 ;
        RECT 53.400 0.310 53.720 0.325 ;
        RECT 51.405 0.080 53.720 0.310 ;
        RECT 51.405 -0.095 51.735 0.080 ;
        RECT 53.400 0.065 53.720 0.080 ;
        RECT 51.460 -0.325 51.690 -0.095 ;
        RECT 51.030 -1.915 52.030 -0.325 ;
        RECT 51.280 -2.545 51.520 -1.915 ;
        RECT 49.110 -2.555 51.520 -2.545 ;
        RECT 48.640 -2.745 51.520 -2.555 ;
        RECT 48.640 -2.785 50.200 -2.745 ;
        RECT 47.690 -3.065 49.590 -3.055 ;
        RECT 47.680 -3.315 49.590 -3.065 ;
        RECT 47.680 -5.485 47.910 -3.315 ;
        RECT 49.070 -3.685 49.300 -3.585 ;
        RECT 51.280 -3.685 51.520 -2.745 ;
        RECT 49.070 -3.925 51.520 -3.685 ;
        RECT 49.070 -4.375 49.300 -3.925 ;
        RECT 49.540 -5.005 49.770 -4.425 ;
        RECT 49.540 -5.135 50.730 -5.005 ;
        RECT 53.960 -5.130 54.230 1.555 ;
        RECT 55.170 -1.585 55.440 1.555 ;
        RECT 55.830 0.310 56.090 0.355 ;
        RECT 57.660 0.310 58.660 0.595 ;
        RECT 61.960 0.310 62.280 0.325 ;
        RECT 55.830 0.080 62.280 0.310 ;
        RECT 55.830 0.035 56.090 0.080 ;
        RECT 57.660 -0.135 58.660 0.080 ;
        RECT 61.960 0.065 62.280 0.080 ;
        RECT 56.780 -0.455 57.100 -0.445 ;
        RECT 57.350 -0.455 59.080 -0.135 ;
        RECT 56.780 -0.695 59.080 -0.455 ;
        RECT 56.780 -0.705 57.100 -0.695 ;
        RECT 57.350 -1.015 59.080 -0.695 ;
        RECT 58.035 -1.365 58.325 -1.315 ;
        RECT 56.550 -1.515 58.325 -1.365 ;
        RECT 54.890 -1.945 55.890 -1.585 ;
        RECT 56.560 -1.945 56.750 -1.515 ;
        RECT 58.035 -1.545 58.325 -1.515 ;
        RECT 62.770 -1.535 63.040 1.555 ;
        RECT 63.520 0.310 63.780 0.355 ;
        RECT 65.250 0.310 66.250 0.645 ;
        RECT 69.780 0.310 70.100 0.325 ;
        RECT 63.520 0.080 70.100 0.310 ;
        RECT 63.520 0.035 63.780 0.080 ;
        RECT 65.250 -0.085 66.250 0.080 ;
        RECT 69.780 0.065 70.100 0.080 ;
        RECT 64.370 -0.405 64.690 -0.395 ;
        RECT 64.940 -0.405 66.670 -0.085 ;
        RECT 64.370 -0.645 66.670 -0.405 ;
        RECT 64.370 -0.655 64.690 -0.645 ;
        RECT 64.940 -0.965 66.670 -0.645 ;
        RECT 65.625 -1.315 65.915 -1.265 ;
        RECT 64.140 -1.465 65.915 -1.315 ;
        RECT 54.890 -2.215 56.750 -1.945 ;
        RECT 54.890 -2.585 55.890 -2.215 ;
        RECT 56.560 -2.715 56.750 -2.215 ;
        RECT 57.080 -1.965 57.340 -1.925 ;
        RECT 57.830 -1.965 58.060 -1.750 ;
        RECT 57.080 -2.205 58.060 -1.965 ;
        RECT 57.080 -2.245 57.340 -2.205 ;
        RECT 57.830 -2.470 58.060 -2.205 ;
        RECT 58.300 -1.805 58.530 -1.750 ;
        RECT 58.730 -1.805 59.050 -1.760 ;
        RECT 58.300 -1.975 59.050 -1.805 ;
        RECT 58.300 -2.470 58.530 -1.975 ;
        RECT 58.730 -2.020 59.050 -1.975 ;
        RECT 62.480 -1.895 63.480 -1.535 ;
        RECT 64.150 -1.895 64.340 -1.465 ;
        RECT 65.625 -1.495 65.915 -1.465 ;
        RECT 70.420 -1.515 70.690 1.555 ;
        RECT 70.960 0.310 71.220 0.355 ;
        RECT 72.860 0.310 73.860 0.665 ;
        RECT 77.760 0.310 78.020 0.355 ;
        RECT 70.960 0.080 78.020 0.310 ;
        RECT 70.960 0.035 71.220 0.080 ;
        RECT 72.860 -0.065 73.860 0.080 ;
        RECT 77.760 0.035 78.020 0.080 ;
        RECT 71.980 -0.385 72.300 -0.375 ;
        RECT 72.550 -0.385 74.280 -0.065 ;
        RECT 71.980 -0.625 74.280 -0.385 ;
        RECT 71.980 -0.635 72.300 -0.625 ;
        RECT 72.550 -0.945 74.280 -0.625 ;
        RECT 73.235 -1.295 73.525 -1.245 ;
        RECT 71.750 -1.445 73.525 -1.295 ;
        RECT 62.480 -2.165 64.340 -1.895 ;
        RECT 62.480 -2.535 63.480 -2.165 ;
        RECT 64.150 -2.665 64.340 -2.165 ;
        RECT 64.670 -1.915 64.930 -1.875 ;
        RECT 65.420 -1.915 65.650 -1.700 ;
        RECT 64.670 -2.155 65.650 -1.915 ;
        RECT 64.670 -2.195 64.930 -2.155 ;
        RECT 65.420 -2.420 65.650 -2.155 ;
        RECT 65.890 -1.755 66.120 -1.700 ;
        RECT 66.320 -1.755 66.640 -1.710 ;
        RECT 65.890 -1.925 66.640 -1.755 ;
        RECT 65.890 -2.420 66.120 -1.925 ;
        RECT 66.320 -1.970 66.640 -1.925 ;
        RECT 70.090 -1.875 71.090 -1.515 ;
        RECT 71.760 -1.875 71.950 -1.445 ;
        RECT 73.235 -1.475 73.525 -1.445 ;
        RECT 78.260 -1.555 78.530 1.555 ;
        RECT 78.880 0.310 79.140 0.355 ;
        RECT 80.860 0.310 81.860 0.625 ;
        RECT 85.370 0.310 85.690 0.325 ;
        RECT 78.880 0.080 85.690 0.310 ;
        RECT 78.880 0.035 79.140 0.080 ;
        RECT 80.860 -0.105 81.860 0.080 ;
        RECT 85.370 0.065 85.690 0.080 ;
        RECT 79.980 -0.425 80.300 -0.415 ;
        RECT 80.550 -0.425 82.280 -0.105 ;
        RECT 79.980 -0.665 82.280 -0.425 ;
        RECT 79.980 -0.675 80.300 -0.665 ;
        RECT 80.550 -0.985 82.280 -0.665 ;
        RECT 81.235 -1.335 81.525 -1.285 ;
        RECT 79.750 -1.485 81.525 -1.335 ;
        RECT 70.090 -2.145 71.950 -1.875 ;
        RECT 70.090 -2.515 71.090 -2.145 ;
        RECT 70.420 -2.575 70.690 -2.515 ;
        RECT 65.625 -2.665 65.915 -2.625 ;
        RECT 71.760 -2.645 71.950 -2.145 ;
        RECT 72.280 -1.895 72.540 -1.855 ;
        RECT 73.030 -1.895 73.260 -1.680 ;
        RECT 72.280 -2.135 73.260 -1.895 ;
        RECT 72.280 -2.175 72.540 -2.135 ;
        RECT 73.030 -2.400 73.260 -2.135 ;
        RECT 73.500 -1.735 73.730 -1.680 ;
        RECT 73.930 -1.735 74.250 -1.690 ;
        RECT 73.500 -1.905 74.250 -1.735 ;
        RECT 73.500 -2.400 73.730 -1.905 ;
        RECT 73.930 -1.950 74.250 -1.905 ;
        RECT 78.090 -1.915 79.090 -1.555 ;
        RECT 79.760 -1.915 79.950 -1.485 ;
        RECT 81.235 -1.515 81.525 -1.485 ;
        RECT 86.180 -1.535 86.450 1.555 ;
        RECT 86.750 0.310 87.010 0.355 ;
        RECT 88.670 0.310 89.670 0.645 ;
        RECT 93.300 0.310 93.620 0.325 ;
        RECT 86.750 0.080 93.620 0.310 ;
        RECT 86.750 0.035 87.010 0.080 ;
        RECT 88.670 -0.085 89.670 0.080 ;
        RECT 93.300 0.065 93.620 0.080 ;
        RECT 87.790 -0.405 88.110 -0.395 ;
        RECT 88.360 -0.405 90.090 -0.085 ;
        RECT 87.790 -0.645 90.090 -0.405 ;
        RECT 87.790 -0.655 88.110 -0.645 ;
        RECT 88.360 -0.965 90.090 -0.645 ;
        RECT 89.045 -1.315 89.335 -1.265 ;
        RECT 87.560 -1.465 89.335 -1.315 ;
        RECT 78.090 -2.185 79.950 -1.915 ;
        RECT 78.090 -2.555 79.090 -2.185 ;
        RECT 73.235 -2.645 73.525 -2.605 ;
        RECT 58.035 -2.715 58.325 -2.675 ;
        RECT 56.560 -2.865 58.350 -2.715 ;
        RECT 64.150 -2.815 65.940 -2.665 ;
        RECT 71.760 -2.795 73.550 -2.645 ;
        RECT 79.760 -2.685 79.950 -2.185 ;
        RECT 80.280 -1.935 80.540 -1.895 ;
        RECT 81.030 -1.935 81.260 -1.720 ;
        RECT 80.280 -2.175 81.260 -1.935 ;
        RECT 80.280 -2.215 80.540 -2.175 ;
        RECT 81.030 -2.440 81.260 -2.175 ;
        RECT 81.500 -1.775 81.730 -1.720 ;
        RECT 81.930 -1.775 82.250 -1.730 ;
        RECT 81.500 -1.945 82.250 -1.775 ;
        RECT 81.500 -2.440 81.730 -1.945 ;
        RECT 81.930 -1.990 82.250 -1.945 ;
        RECT 85.900 -1.895 86.900 -1.535 ;
        RECT 87.570 -1.895 87.760 -1.465 ;
        RECT 89.045 -1.495 89.335 -1.465 ;
        RECT 93.850 -1.555 94.120 1.555 ;
        RECT 94.510 0.310 94.770 0.355 ;
        RECT 96.260 0.310 97.260 0.625 ;
        RECT 100.530 0.310 100.850 0.325 ;
        RECT 94.510 0.080 100.850 0.310 ;
        RECT 94.510 0.035 94.770 0.080 ;
        RECT 96.260 -0.105 97.260 0.080 ;
        RECT 100.530 0.065 100.850 0.080 ;
        RECT 95.380 -0.425 95.700 -0.415 ;
        RECT 95.950 -0.425 97.680 -0.105 ;
        RECT 95.380 -0.665 97.680 -0.425 ;
        RECT 95.380 -0.675 95.700 -0.665 ;
        RECT 95.950 -0.985 97.680 -0.665 ;
        RECT 96.635 -1.335 96.925 -1.285 ;
        RECT 95.150 -1.485 96.925 -1.335 ;
        RECT 85.900 -2.165 87.760 -1.895 ;
        RECT 85.900 -2.535 86.900 -2.165 ;
        RECT 86.180 -2.575 86.450 -2.535 ;
        RECT 81.235 -2.685 81.525 -2.645 ;
        RECT 87.570 -2.665 87.760 -2.165 ;
        RECT 88.090 -1.915 88.350 -1.875 ;
        RECT 88.840 -1.915 89.070 -1.700 ;
        RECT 88.090 -2.155 89.070 -1.915 ;
        RECT 88.090 -2.195 88.350 -2.155 ;
        RECT 88.840 -2.420 89.070 -2.155 ;
        RECT 89.310 -1.755 89.540 -1.700 ;
        RECT 89.740 -1.755 90.060 -1.710 ;
        RECT 89.310 -1.925 90.060 -1.755 ;
        RECT 89.310 -2.420 89.540 -1.925 ;
        RECT 89.740 -1.970 90.060 -1.925 ;
        RECT 93.490 -1.915 94.490 -1.555 ;
        RECT 95.160 -1.915 95.350 -1.485 ;
        RECT 96.635 -1.515 96.925 -1.485 ;
        RECT 101.150 -1.585 101.420 1.555 ;
        RECT 102.685 1.475 102.975 2.655 ;
        RECT 107.130 1.710 107.470 3.920 ;
        RECT 114.380 4.125 118.270 4.345 ;
        RECT 114.380 4.110 116.330 4.125 ;
        RECT 112.560 1.475 113.140 3.370 ;
        RECT 102.685 1.185 113.140 1.475 ;
        RECT 101.610 0.310 101.870 0.355 ;
        RECT 103.650 0.310 104.650 0.595 ;
        RECT 107.100 0.570 107.500 0.910 ;
        RECT 101.610 0.305 104.650 0.310 ;
        RECT 107.130 0.305 107.470 0.570 ;
        RECT 101.610 0.080 110.715 0.305 ;
        RECT 101.610 0.035 101.870 0.080 ;
        RECT 103.650 0.055 110.715 0.080 ;
        RECT 103.650 -0.135 104.650 0.055 ;
        RECT 102.770 -0.455 103.090 -0.445 ;
        RECT 103.340 -0.455 105.070 -0.135 ;
        RECT 102.770 -0.695 105.070 -0.455 ;
        RECT 102.770 -0.705 103.090 -0.695 ;
        RECT 103.340 -1.015 105.070 -0.695 ;
        RECT 104.025 -1.365 104.315 -1.315 ;
        RECT 102.540 -1.515 104.315 -1.365 ;
        RECT 93.490 -2.185 95.350 -1.915 ;
        RECT 93.490 -2.555 94.490 -2.185 ;
        RECT 93.850 -2.565 94.120 -2.555 ;
        RECT 89.045 -2.665 89.335 -2.625 ;
        RECT 65.625 -2.855 65.915 -2.815 ;
        RECT 73.235 -2.835 73.525 -2.795 ;
        RECT 79.760 -2.835 81.550 -2.685 ;
        RECT 87.570 -2.815 89.360 -2.665 ;
        RECT 95.160 -2.685 95.350 -2.185 ;
        RECT 95.680 -1.935 95.940 -1.895 ;
        RECT 96.430 -1.935 96.660 -1.720 ;
        RECT 95.680 -2.175 96.660 -1.935 ;
        RECT 95.680 -2.215 95.940 -2.175 ;
        RECT 96.430 -2.440 96.660 -2.175 ;
        RECT 96.900 -1.775 97.130 -1.720 ;
        RECT 97.330 -1.775 97.650 -1.730 ;
        RECT 96.900 -1.945 97.650 -1.775 ;
        RECT 96.900 -2.440 97.130 -1.945 ;
        RECT 97.330 -1.990 97.650 -1.945 ;
        RECT 100.880 -1.945 101.880 -1.585 ;
        RECT 102.550 -1.945 102.740 -1.515 ;
        RECT 104.025 -1.545 104.315 -1.515 ;
        RECT 110.465 -1.635 110.715 0.055 ;
        RECT 100.880 -2.215 102.740 -1.945 ;
        RECT 100.880 -2.585 101.880 -2.215 ;
        RECT 96.635 -2.685 96.925 -2.645 ;
        RECT 58.035 -2.905 58.325 -2.865 ;
        RECT 81.235 -2.875 81.525 -2.835 ;
        RECT 89.045 -2.855 89.335 -2.815 ;
        RECT 95.160 -2.835 96.950 -2.685 ;
        RECT 102.550 -2.715 102.740 -2.215 ;
        RECT 103.070 -1.965 103.330 -1.925 ;
        RECT 103.820 -1.965 104.050 -1.750 ;
        RECT 103.070 -2.205 104.050 -1.965 ;
        RECT 103.070 -2.245 103.330 -2.205 ;
        RECT 103.820 -2.470 104.050 -2.205 ;
        RECT 104.290 -1.805 104.520 -1.750 ;
        RECT 104.720 -1.805 105.040 -1.760 ;
        RECT 104.290 -1.975 105.040 -1.805 ;
        RECT 104.290 -2.470 104.520 -1.975 ;
        RECT 104.720 -2.020 105.040 -1.975 ;
        RECT 110.190 -2.365 111.190 -1.635 ;
        RECT 109.310 -2.645 109.630 -2.605 ;
        RECT 109.830 -2.645 111.560 -2.365 ;
        RECT 104.025 -2.715 104.315 -2.675 ;
        RECT 96.635 -2.875 96.925 -2.835 ;
        RECT 102.550 -2.865 104.340 -2.715 ;
        RECT 109.310 -2.825 111.560 -2.645 ;
        RECT 109.310 -2.865 109.630 -2.825 ;
        RECT 104.025 -2.905 104.315 -2.865 ;
        RECT 109.830 -3.135 111.560 -2.825 ;
        RECT 110.545 -3.475 110.835 -3.445 ;
        RECT 108.710 -3.665 110.850 -3.475 ;
        RECT 73.235 -4.075 73.525 -4.065 ;
        RECT 108.720 -4.075 108.900 -3.665 ;
        RECT 110.545 -3.675 110.835 -3.665 ;
        RECT 65.625 -4.095 65.915 -4.085 ;
        RECT 58.035 -4.145 58.325 -4.135 ;
        RECT 55.850 -4.385 58.330 -4.145 ;
        RECT 63.440 -4.335 65.920 -4.095 ;
        RECT 71.050 -4.315 73.530 -4.075 ;
        RECT 89.045 -4.095 89.335 -4.085 ;
        RECT 81.235 -4.115 81.525 -4.105 ;
        RECT 55.880 -4.825 56.100 -4.385 ;
        RECT 51.190 -5.135 54.230 -5.130 ;
        RECT 49.540 -5.205 54.230 -5.135 ;
        RECT 49.540 -5.215 49.770 -5.205 ;
        RECT 50.490 -5.400 54.230 -5.205 ;
        RECT 55.450 -5.105 56.110 -4.825 ;
        RECT 57.370 -4.845 57.690 -4.785 ;
        RECT 57.830 -4.845 58.060 -4.570 ;
        RECT 57.370 -4.985 58.060 -4.845 ;
        RECT 57.370 -5.045 57.690 -4.985 ;
        RECT 47.680 -5.745 49.590 -5.485 ;
        RECT 47.680 -6.630 47.910 -5.745 ;
        RECT 50.490 -6.630 50.700 -5.400 ;
        RECT 47.680 -6.860 50.700 -6.630 ;
        RECT 48.420 -7.190 48.740 -7.165 ;
        RECT 50.490 -7.190 50.700 -6.860 ;
        RECT 54.250 -6.205 55.250 -5.905 ;
        RECT 55.450 -6.205 55.730 -5.105 ;
        RECT 55.880 -5.505 56.100 -5.105 ;
        RECT 57.830 -5.290 58.060 -4.985 ;
        RECT 58.300 -5.075 58.530 -4.570 ;
        RECT 63.470 -4.775 63.690 -4.335 ;
        RECT 63.040 -5.055 63.700 -4.775 ;
        RECT 64.960 -4.795 65.280 -4.735 ;
        RECT 65.420 -4.795 65.650 -4.520 ;
        RECT 64.960 -4.935 65.650 -4.795 ;
        RECT 64.960 -4.995 65.280 -4.935 ;
        RECT 59.300 -5.075 59.480 -5.070 ;
        RECT 58.300 -5.245 59.490 -5.075 ;
        RECT 58.300 -5.290 58.530 -5.245 ;
        RECT 58.035 -5.505 58.325 -5.495 ;
        RECT 55.880 -5.745 58.360 -5.505 ;
        RECT 59.300 -6.035 59.480 -5.245 ;
        RECT 60.140 -6.035 61.140 -5.635 ;
        RECT 54.250 -6.485 55.730 -6.205 ;
        RECT 59.290 -6.055 61.140 -6.035 ;
        RECT 61.840 -6.055 62.840 -5.855 ;
        RECT 59.290 -6.155 62.840 -6.055 ;
        RECT 63.040 -6.155 63.320 -5.055 ;
        RECT 63.470 -5.455 63.690 -5.055 ;
        RECT 65.420 -5.240 65.650 -4.935 ;
        RECT 65.890 -5.025 66.120 -4.520 ;
        RECT 71.080 -4.755 71.300 -4.315 ;
        RECT 79.050 -4.355 81.530 -4.115 ;
        RECT 86.860 -4.335 89.340 -4.095 ;
        RECT 96.635 -4.115 96.925 -4.105 ;
        RECT 66.890 -5.025 67.070 -5.020 ;
        RECT 65.890 -5.195 67.080 -5.025 ;
        RECT 70.650 -5.035 71.310 -4.755 ;
        RECT 72.570 -4.775 72.890 -4.715 ;
        RECT 73.030 -4.775 73.260 -4.500 ;
        RECT 72.570 -4.915 73.260 -4.775 ;
        RECT 72.570 -4.975 72.890 -4.915 ;
        RECT 65.890 -5.240 66.120 -5.195 ;
        RECT 65.625 -5.455 65.915 -5.445 ;
        RECT 63.470 -5.695 65.950 -5.455 ;
        RECT 66.890 -5.985 67.070 -5.195 ;
        RECT 67.730 -5.915 68.730 -5.585 ;
        RECT 69.450 -5.915 70.450 -5.835 ;
        RECT 67.730 -5.985 70.450 -5.915 ;
        RECT 59.290 -6.255 63.320 -6.155 ;
        RECT 66.880 -6.135 70.450 -5.985 ;
        RECT 70.650 -6.135 70.930 -5.035 ;
        RECT 71.080 -5.435 71.300 -5.035 ;
        RECT 73.030 -5.220 73.260 -4.915 ;
        RECT 73.500 -5.005 73.730 -4.500 ;
        RECT 79.080 -4.795 79.300 -4.355 ;
        RECT 74.500 -5.005 74.680 -5.000 ;
        RECT 73.500 -5.175 74.690 -5.005 ;
        RECT 78.650 -5.075 79.310 -4.795 ;
        RECT 80.570 -4.815 80.890 -4.755 ;
        RECT 81.030 -4.815 81.260 -4.540 ;
        RECT 80.570 -4.955 81.260 -4.815 ;
        RECT 80.570 -5.015 80.890 -4.955 ;
        RECT 73.500 -5.220 73.730 -5.175 ;
        RECT 73.235 -5.435 73.525 -5.425 ;
        RECT 71.080 -5.675 73.560 -5.435 ;
        RECT 74.500 -5.965 74.680 -5.175 ;
        RECT 75.340 -5.915 76.340 -5.565 ;
        RECT 77.450 -5.915 78.450 -5.875 ;
        RECT 75.340 -5.965 78.450 -5.915 ;
        RECT 66.880 -6.205 70.930 -6.135 ;
        RECT 74.490 -6.175 78.450 -5.965 ;
        RECT 78.650 -6.175 78.930 -5.075 ;
        RECT 79.080 -5.475 79.300 -5.075 ;
        RECT 81.030 -5.260 81.260 -4.955 ;
        RECT 81.500 -5.045 81.730 -4.540 ;
        RECT 86.890 -4.775 87.110 -4.335 ;
        RECT 94.450 -4.355 96.930 -4.115 ;
        RECT 104.025 -4.145 104.315 -4.135 ;
        RECT 82.500 -5.045 82.680 -5.040 ;
        RECT 81.500 -5.215 82.690 -5.045 ;
        RECT 86.460 -5.055 87.120 -4.775 ;
        RECT 88.380 -4.795 88.700 -4.735 ;
        RECT 88.840 -4.795 89.070 -4.520 ;
        RECT 88.380 -4.935 89.070 -4.795 ;
        RECT 88.380 -4.995 88.700 -4.935 ;
        RECT 81.500 -5.260 81.730 -5.215 ;
        RECT 81.235 -5.475 81.525 -5.465 ;
        RECT 79.080 -5.715 81.560 -5.475 ;
        RECT 82.500 -6.005 82.680 -5.215 ;
        RECT 83.340 -5.955 84.340 -5.605 ;
        RECT 85.260 -5.955 86.260 -5.855 ;
        RECT 83.340 -6.005 86.260 -5.955 ;
        RECT 74.490 -6.185 78.930 -6.175 ;
        RECT 54.250 -6.905 55.250 -6.485 ;
        RECT 48.420 -7.400 50.700 -7.190 ;
        RECT 48.420 -7.425 48.740 -7.400 ;
        RECT 54.535 -7.620 54.805 -6.905 ;
        RECT 52.625 -7.890 54.805 -7.620 ;
        RECT 55.440 -7.635 55.720 -6.485 ;
        RECT 57.080 -6.755 57.400 -6.715 ;
        RECT 59.300 -6.755 59.480 -6.255 ;
        RECT 60.140 -6.415 63.320 -6.255 ;
        RECT 60.140 -6.635 61.140 -6.415 ;
        RECT 61.840 -6.435 63.320 -6.415 ;
        RECT 57.080 -6.935 59.480 -6.755 ;
        RECT 61.840 -6.855 62.840 -6.435 ;
        RECT 57.080 -6.975 57.400 -6.935 ;
        RECT 59.300 -6.955 59.480 -6.935 ;
        RECT 55.880 -7.505 58.360 -7.265 ;
        RECT 55.880 -7.635 56.070 -7.505 ;
        RECT 58.045 -7.515 58.335 -7.505 ;
        RECT 44.410 -8.555 45.410 -8.135 ;
        RECT 47.730 -8.145 49.570 -7.915 ;
        RECT 47.750 -8.460 47.950 -8.145 ;
        RECT 49.265 -8.155 49.555 -8.145 ;
        RECT 47.215 -8.555 47.950 -8.460 ;
        RECT 44.410 -8.730 47.950 -8.555 ;
        RECT 48.420 -8.400 48.740 -8.375 ;
        RECT 49.060 -8.400 49.290 -8.315 ;
        RECT 48.420 -8.610 49.290 -8.400 ;
        RECT 48.420 -8.635 48.740 -8.610 ;
        RECT 44.410 -8.825 47.485 -8.730 ;
        RECT 44.410 -9.135 45.410 -8.825 ;
        RECT 40.950 -10.940 46.840 -10.600 ;
        RECT 18.390 -11.640 18.590 -11.610 ;
        RECT 33.185 -11.615 33.450 -11.375 ;
        RECT 17.690 -11.710 17.880 -11.665 ;
        RECT 18.145 -11.870 24.215 -11.640 ;
        RECT 33.220 -11.665 33.450 -11.615 ;
        RECT 17.120 -12.740 17.320 -12.380 ;
        RECT 18.390 -12.740 18.590 -11.870 ;
        RECT 17.120 -12.940 18.590 -12.740 ;
        RECT 40.950 -14.290 41.390 -10.940 ;
        RECT 47.215 -13.175 47.485 -8.825 ;
        RECT 47.750 -8.885 47.950 -8.730 ;
        RECT 49.060 -8.735 49.290 -8.610 ;
        RECT 49.530 -8.465 49.760 -8.315 ;
        RECT 49.530 -8.685 50.780 -8.465 ;
        RECT 49.530 -8.735 49.760 -8.685 ;
        RECT 47.740 -9.115 49.580 -8.885 ;
        RECT 49.265 -9.125 49.555 -9.115 ;
        RECT 48.630 -9.485 50.190 -9.405 ;
        RECT 48.600 -9.775 50.210 -9.485 ;
        RECT 50.560 -9.775 50.780 -8.685 ;
        RECT 48.600 -9.995 50.780 -9.775 ;
        RECT 48.600 -10.355 50.210 -9.995 ;
        RECT 48.080 -10.600 48.420 -10.570 ;
        RECT 48.880 -10.600 49.880 -10.355 ;
        RECT 48.080 -10.940 49.880 -10.600 ;
        RECT 48.080 -10.970 48.420 -10.940 ;
        RECT 48.880 -10.985 49.880 -10.940 ;
        RECT 49.460 -11.965 49.700 -10.985 ;
        RECT 52.050 -11.965 52.370 -11.955 ;
        RECT 49.460 -12.205 52.370 -11.965 ;
        RECT 52.050 -12.215 52.370 -12.205 ;
        RECT 51.125 -13.175 51.395 -13.145 ;
        RECT 47.215 -13.445 51.395 -13.175 ;
        RECT 51.125 -13.475 51.395 -13.445 ;
        RECT 52.625 -13.930 52.895 -7.890 ;
        RECT 55.440 -7.915 56.070 -7.635 ;
        RECT 63.030 -7.585 63.310 -6.435 ;
        RECT 64.670 -6.705 64.990 -6.665 ;
        RECT 66.890 -6.705 67.070 -6.205 ;
        RECT 67.730 -6.275 70.930 -6.205 ;
        RECT 67.730 -6.585 68.730 -6.275 ;
        RECT 69.450 -6.415 70.930 -6.275 ;
        RECT 64.670 -6.885 67.070 -6.705 ;
        RECT 69.450 -6.835 70.450 -6.415 ;
        RECT 64.670 -6.925 64.990 -6.885 ;
        RECT 66.890 -6.905 67.070 -6.885 ;
        RECT 63.470 -7.455 65.950 -7.215 ;
        RECT 63.470 -7.585 63.660 -7.455 ;
        RECT 65.635 -7.465 65.925 -7.455 ;
        RECT 55.880 -8.245 56.070 -7.915 ;
        RECT 57.110 -7.745 57.370 -7.675 ;
        RECT 57.840 -7.745 58.070 -7.675 ;
        RECT 57.110 -7.925 58.070 -7.745 ;
        RECT 57.110 -7.995 57.370 -7.925 ;
        RECT 57.690 -7.935 58.070 -7.925 ;
        RECT 57.840 -8.095 58.070 -7.935 ;
        RECT 58.310 -7.865 58.540 -7.675 ;
        RECT 63.030 -7.865 63.660 -7.585 ;
        RECT 70.640 -7.565 70.920 -6.415 ;
        RECT 72.280 -6.685 72.600 -6.645 ;
        RECT 74.500 -6.685 74.680 -6.185 ;
        RECT 75.340 -6.275 78.930 -6.185 ;
        RECT 82.490 -6.155 86.260 -6.005 ;
        RECT 86.460 -6.155 86.740 -5.055 ;
        RECT 86.890 -5.455 87.110 -5.055 ;
        RECT 88.840 -5.240 89.070 -4.935 ;
        RECT 89.310 -5.025 89.540 -4.520 ;
        RECT 94.480 -4.795 94.700 -4.355 ;
        RECT 101.840 -4.385 104.320 -4.145 ;
        RECT 108.120 -4.325 108.900 -4.075 ;
        RECT 90.310 -5.025 90.490 -5.020 ;
        RECT 89.310 -5.195 90.500 -5.025 ;
        RECT 94.050 -5.075 94.710 -4.795 ;
        RECT 95.970 -4.815 96.290 -4.755 ;
        RECT 96.430 -4.815 96.660 -4.540 ;
        RECT 95.970 -4.955 96.660 -4.815 ;
        RECT 95.970 -5.015 96.290 -4.955 ;
        RECT 89.310 -5.240 89.540 -5.195 ;
        RECT 89.045 -5.455 89.335 -5.445 ;
        RECT 86.890 -5.695 89.370 -5.455 ;
        RECT 90.310 -5.985 90.490 -5.195 ;
        RECT 91.150 -5.955 92.150 -5.585 ;
        RECT 92.850 -5.955 93.850 -5.875 ;
        RECT 91.150 -5.985 93.850 -5.955 ;
        RECT 82.490 -6.225 86.740 -6.155 ;
        RECT 90.300 -6.175 93.850 -5.985 ;
        RECT 94.050 -6.175 94.330 -5.075 ;
        RECT 94.480 -5.475 94.700 -5.075 ;
        RECT 96.430 -5.260 96.660 -4.955 ;
        RECT 96.900 -5.045 97.130 -4.540 ;
        RECT 101.870 -4.825 102.090 -4.385 ;
        RECT 97.900 -5.045 98.080 -5.040 ;
        RECT 96.900 -5.215 98.090 -5.045 ;
        RECT 101.440 -5.105 102.100 -4.825 ;
        RECT 103.360 -4.845 103.680 -4.785 ;
        RECT 103.820 -4.845 104.050 -4.570 ;
        RECT 103.360 -4.985 104.050 -4.845 ;
        RECT 103.360 -5.045 103.680 -4.985 ;
        RECT 96.900 -5.260 97.130 -5.215 ;
        RECT 96.635 -5.475 96.925 -5.465 ;
        RECT 94.480 -5.715 96.960 -5.475 ;
        RECT 97.900 -6.005 98.080 -5.215 ;
        RECT 98.740 -6.005 99.740 -5.605 ;
        RECT 100.240 -6.005 101.240 -5.905 ;
        RECT 90.300 -6.205 94.330 -6.175 ;
        RECT 75.340 -6.565 76.340 -6.275 ;
        RECT 77.450 -6.455 78.930 -6.275 ;
        RECT 72.280 -6.865 74.680 -6.685 ;
        RECT 72.280 -6.905 72.600 -6.865 ;
        RECT 74.500 -6.885 74.680 -6.865 ;
        RECT 77.450 -6.875 78.450 -6.455 ;
        RECT 71.080 -7.435 73.560 -7.195 ;
        RECT 71.080 -7.565 71.270 -7.435 ;
        RECT 73.245 -7.445 73.535 -7.435 ;
        RECT 58.310 -8.035 59.490 -7.865 ;
        RECT 58.310 -8.095 58.540 -8.035 ;
        RECT 55.880 -8.485 58.360 -8.245 ;
        RECT 57.180 -9.390 57.500 -9.345 ;
        RECT 59.315 -9.390 59.485 -8.035 ;
        RECT 63.470 -8.195 63.660 -7.865 ;
        RECT 64.700 -7.695 64.960 -7.625 ;
        RECT 65.430 -7.695 65.660 -7.625 ;
        RECT 64.700 -7.875 65.660 -7.695 ;
        RECT 64.700 -7.945 64.960 -7.875 ;
        RECT 65.280 -7.885 65.660 -7.875 ;
        RECT 65.430 -8.045 65.660 -7.885 ;
        RECT 65.900 -7.815 66.130 -7.625 ;
        RECT 65.900 -7.985 67.080 -7.815 ;
        RECT 70.640 -7.845 71.270 -7.565 ;
        RECT 78.640 -7.605 78.920 -6.455 ;
        RECT 80.280 -6.725 80.600 -6.685 ;
        RECT 82.500 -6.725 82.680 -6.225 ;
        RECT 83.340 -6.315 86.740 -6.225 ;
        RECT 83.340 -6.605 84.340 -6.315 ;
        RECT 85.260 -6.435 86.740 -6.315 ;
        RECT 80.280 -6.905 82.680 -6.725 ;
        RECT 85.260 -6.855 86.260 -6.435 ;
        RECT 80.280 -6.945 80.600 -6.905 ;
        RECT 82.500 -6.925 82.680 -6.905 ;
        RECT 79.080 -7.475 81.560 -7.235 ;
        RECT 79.080 -7.605 79.270 -7.475 ;
        RECT 81.245 -7.485 81.535 -7.475 ;
        RECT 65.900 -8.045 66.130 -7.985 ;
        RECT 63.470 -8.435 65.950 -8.195 ;
        RECT 57.180 -9.560 59.485 -9.390 ;
        RECT 64.770 -9.340 65.090 -9.295 ;
        RECT 66.905 -9.340 67.075 -7.985 ;
        RECT 71.080 -8.175 71.270 -7.845 ;
        RECT 72.310 -7.675 72.570 -7.605 ;
        RECT 73.040 -7.675 73.270 -7.605 ;
        RECT 72.310 -7.855 73.270 -7.675 ;
        RECT 72.310 -7.925 72.570 -7.855 ;
        RECT 72.890 -7.865 73.270 -7.855 ;
        RECT 73.040 -8.025 73.270 -7.865 ;
        RECT 73.510 -7.795 73.740 -7.605 ;
        RECT 73.510 -7.965 74.690 -7.795 ;
        RECT 78.640 -7.885 79.270 -7.605 ;
        RECT 86.450 -7.585 86.730 -6.435 ;
        RECT 88.090 -6.705 88.410 -6.665 ;
        RECT 90.310 -6.705 90.490 -6.205 ;
        RECT 91.150 -6.315 94.330 -6.205 ;
        RECT 97.890 -6.205 101.240 -6.005 ;
        RECT 101.440 -6.205 101.720 -5.105 ;
        RECT 101.870 -5.505 102.090 -5.105 ;
        RECT 103.820 -5.290 104.050 -4.985 ;
        RECT 104.290 -5.075 104.520 -4.570 ;
        RECT 105.290 -5.075 105.470 -5.070 ;
        RECT 104.290 -5.245 105.480 -5.075 ;
        RECT 104.290 -5.290 104.520 -5.245 ;
        RECT 104.025 -5.505 104.315 -5.495 ;
        RECT 101.870 -5.745 104.350 -5.505 ;
        RECT 105.290 -6.035 105.470 -5.245 ;
        RECT 106.130 -5.955 107.130 -5.635 ;
        RECT 108.130 -5.955 108.300 -4.325 ;
        RECT 108.720 -4.815 108.900 -4.325 ;
        RECT 109.340 -4.125 109.600 -4.055 ;
        RECT 110.340 -4.125 110.570 -3.880 ;
        RECT 109.340 -4.305 110.570 -4.125 ;
        RECT 109.340 -4.375 109.600 -4.305 ;
        RECT 110.340 -4.600 110.570 -4.305 ;
        RECT 110.810 -4.135 111.040 -3.880 ;
        RECT 110.810 -4.325 112.010 -4.135 ;
        RECT 110.810 -4.600 111.040 -4.325 ;
        RECT 110.545 -4.815 110.835 -4.805 ;
        RECT 108.720 -5.005 110.860 -4.815 ;
        RECT 110.545 -5.035 110.835 -5.005 ;
        RECT 106.130 -6.035 108.300 -5.955 ;
        RECT 97.890 -6.225 101.720 -6.205 ;
        RECT 91.150 -6.585 92.150 -6.315 ;
        RECT 92.850 -6.455 94.330 -6.315 ;
        RECT 88.090 -6.885 90.490 -6.705 ;
        RECT 92.850 -6.875 93.850 -6.455 ;
        RECT 88.090 -6.925 88.410 -6.885 ;
        RECT 90.310 -6.905 90.490 -6.885 ;
        RECT 86.890 -7.455 89.370 -7.215 ;
        RECT 86.890 -7.585 87.080 -7.455 ;
        RECT 89.055 -7.465 89.345 -7.455 ;
        RECT 73.510 -8.025 73.740 -7.965 ;
        RECT 71.080 -8.415 73.560 -8.175 ;
        RECT 64.770 -9.510 67.075 -9.340 ;
        RECT 72.380 -9.320 72.700 -9.275 ;
        RECT 74.515 -9.320 74.685 -7.965 ;
        RECT 79.080 -8.215 79.270 -7.885 ;
        RECT 80.310 -7.715 80.570 -7.645 ;
        RECT 81.040 -7.715 81.270 -7.645 ;
        RECT 80.310 -7.895 81.270 -7.715 ;
        RECT 80.310 -7.965 80.570 -7.895 ;
        RECT 80.890 -7.905 81.270 -7.895 ;
        RECT 81.040 -8.065 81.270 -7.905 ;
        RECT 81.510 -7.835 81.740 -7.645 ;
        RECT 81.510 -8.005 82.690 -7.835 ;
        RECT 86.450 -7.865 87.080 -7.585 ;
        RECT 94.040 -7.605 94.320 -6.455 ;
        RECT 95.680 -6.725 96.000 -6.685 ;
        RECT 97.900 -6.725 98.080 -6.225 ;
        RECT 98.740 -6.365 101.720 -6.225 ;
        RECT 105.280 -6.225 108.300 -6.035 ;
        RECT 111.815 -5.425 112.005 -4.325 ;
        RECT 112.850 -4.935 113.140 1.185 ;
        RECT 112.470 -5.425 113.470 -4.935 ;
        RECT 111.815 -5.685 113.470 -5.425 ;
        RECT 105.280 -6.255 107.130 -6.225 ;
        RECT 98.740 -6.605 99.740 -6.365 ;
        RECT 100.240 -6.485 101.720 -6.365 ;
        RECT 95.680 -6.905 98.080 -6.725 ;
        RECT 100.240 -6.905 101.240 -6.485 ;
        RECT 95.680 -6.945 96.000 -6.905 ;
        RECT 97.900 -6.925 98.080 -6.905 ;
        RECT 94.480 -7.475 96.960 -7.235 ;
        RECT 94.480 -7.605 94.670 -7.475 ;
        RECT 96.645 -7.485 96.935 -7.475 ;
        RECT 81.510 -8.065 81.740 -8.005 ;
        RECT 79.080 -8.455 81.560 -8.215 ;
        RECT 72.380 -9.490 74.685 -9.320 ;
        RECT 80.380 -9.360 80.700 -9.315 ;
        RECT 82.515 -9.360 82.685 -8.005 ;
        RECT 86.890 -8.195 87.080 -7.865 ;
        RECT 88.120 -7.695 88.380 -7.625 ;
        RECT 88.850 -7.695 89.080 -7.625 ;
        RECT 88.120 -7.875 89.080 -7.695 ;
        RECT 88.120 -7.945 88.380 -7.875 ;
        RECT 88.700 -7.885 89.080 -7.875 ;
        RECT 88.850 -8.045 89.080 -7.885 ;
        RECT 89.320 -7.815 89.550 -7.625 ;
        RECT 89.320 -7.985 90.500 -7.815 ;
        RECT 94.040 -7.885 94.670 -7.605 ;
        RECT 101.430 -7.635 101.710 -6.485 ;
        RECT 103.070 -6.755 103.390 -6.715 ;
        RECT 105.290 -6.755 105.470 -6.255 ;
        RECT 106.130 -6.635 107.130 -6.255 ;
        RECT 103.070 -6.935 105.470 -6.755 ;
        RECT 103.070 -6.975 103.390 -6.935 ;
        RECT 105.290 -6.955 105.470 -6.935 ;
        RECT 101.870 -7.505 104.350 -7.265 ;
        RECT 101.870 -7.635 102.060 -7.505 ;
        RECT 104.035 -7.515 104.325 -7.505 ;
        RECT 89.320 -8.045 89.550 -7.985 ;
        RECT 86.890 -8.435 89.370 -8.195 ;
        RECT 64.770 -9.555 65.090 -9.510 ;
        RECT 72.380 -9.535 72.700 -9.490 ;
        RECT 80.380 -9.530 82.685 -9.360 ;
        RECT 88.190 -9.340 88.510 -9.295 ;
        RECT 90.325 -9.340 90.495 -7.985 ;
        RECT 94.480 -8.215 94.670 -7.885 ;
        RECT 95.710 -7.715 95.970 -7.645 ;
        RECT 96.440 -7.715 96.670 -7.645 ;
        RECT 95.710 -7.895 96.670 -7.715 ;
        RECT 95.710 -7.965 95.970 -7.895 ;
        RECT 96.290 -7.905 96.670 -7.895 ;
        RECT 96.440 -8.065 96.670 -7.905 ;
        RECT 96.910 -7.835 97.140 -7.645 ;
        RECT 96.910 -8.005 98.090 -7.835 ;
        RECT 101.430 -7.915 102.060 -7.635 ;
        RECT 96.910 -8.065 97.140 -8.005 ;
        RECT 94.480 -8.455 96.960 -8.215 ;
        RECT 88.190 -9.510 90.495 -9.340 ;
        RECT 95.780 -9.360 96.100 -9.315 ;
        RECT 97.915 -9.360 98.085 -8.005 ;
        RECT 101.870 -8.245 102.060 -7.915 ;
        RECT 103.100 -7.745 103.360 -7.675 ;
        RECT 103.830 -7.745 104.060 -7.675 ;
        RECT 103.100 -7.925 104.060 -7.745 ;
        RECT 103.100 -7.995 103.360 -7.925 ;
        RECT 103.680 -7.935 104.060 -7.925 ;
        RECT 103.830 -8.095 104.060 -7.935 ;
        RECT 104.300 -7.865 104.530 -7.675 ;
        RECT 104.300 -8.035 105.480 -7.865 ;
        RECT 104.300 -8.095 104.530 -8.035 ;
        RECT 101.870 -8.485 104.350 -8.245 ;
        RECT 57.180 -9.605 57.500 -9.560 ;
        RECT 80.380 -9.575 80.700 -9.530 ;
        RECT 88.190 -9.555 88.510 -9.510 ;
        RECT 95.780 -9.530 98.085 -9.360 ;
        RECT 103.170 -9.390 103.490 -9.345 ;
        RECT 105.305 -9.390 105.475 -8.035 ;
        RECT 95.780 -9.575 96.100 -9.530 ;
        RECT 103.170 -9.560 105.475 -9.390 ;
        RECT 103.170 -9.605 103.490 -9.560 ;
        RECT 65.645 -9.695 65.935 -9.665 ;
        RECT 73.255 -9.675 73.545 -9.645 ;
        RECT 58.055 -9.745 58.345 -9.715 ;
        RECT 55.200 -10.035 56.200 -9.805 ;
        RECT 56.500 -9.965 58.360 -9.745 ;
        RECT 56.500 -10.035 56.720 -9.965 ;
        RECT 55.200 -10.255 56.720 -10.035 ;
        RECT 62.790 -9.985 63.790 -9.755 ;
        RECT 64.090 -9.915 65.950 -9.695 ;
        RECT 64.090 -9.985 64.310 -9.915 ;
        RECT 57.180 -10.230 57.500 -10.185 ;
        RECT 57.850 -10.230 58.080 -10.105 ;
        RECT 55.200 -10.805 56.200 -10.255 ;
        RECT 56.490 -10.685 56.710 -10.255 ;
        RECT 57.180 -10.400 58.080 -10.230 ;
        RECT 57.180 -10.445 57.500 -10.400 ;
        RECT 57.760 -10.430 58.080 -10.400 ;
        RECT 57.850 -10.525 58.080 -10.430 ;
        RECT 58.320 -10.285 58.550 -10.105 ;
        RECT 62.790 -10.205 64.310 -9.985 ;
        RECT 70.400 -9.965 71.400 -9.735 ;
        RECT 71.700 -9.895 73.560 -9.675 ;
        RECT 81.255 -9.715 81.545 -9.685 ;
        RECT 89.065 -9.695 89.355 -9.665 ;
        RECT 71.700 -9.965 71.920 -9.895 ;
        RECT 64.770 -10.180 65.090 -10.135 ;
        RECT 65.440 -10.180 65.670 -10.055 ;
        RECT 58.320 -10.455 59.050 -10.285 ;
        RECT 58.320 -10.525 58.550 -10.455 ;
        RECT 53.300 -11.965 53.560 -11.925 ;
        RECT 54.910 -11.965 55.230 -11.955 ;
        RECT 53.300 -12.205 55.230 -11.965 ;
        RECT 53.300 -12.245 53.560 -12.205 ;
        RECT 54.910 -12.215 55.230 -12.205 ;
        RECT 55.450 -13.175 55.720 -10.805 ;
        RECT 56.490 -10.905 58.345 -10.685 ;
        RECT 58.055 -10.915 58.345 -10.905 ;
        RECT 58.855 -11.105 59.025 -10.455 ;
        RECT 62.790 -10.755 63.790 -10.205 ;
        RECT 64.080 -10.635 64.300 -10.205 ;
        RECT 64.770 -10.350 65.670 -10.180 ;
        RECT 64.770 -10.395 65.090 -10.350 ;
        RECT 65.350 -10.380 65.670 -10.350 ;
        RECT 65.440 -10.475 65.670 -10.380 ;
        RECT 65.910 -10.235 66.140 -10.055 ;
        RECT 70.400 -10.185 71.920 -9.965 ;
        RECT 78.400 -10.005 79.400 -9.775 ;
        RECT 79.700 -9.935 81.560 -9.715 ;
        RECT 79.700 -10.005 79.920 -9.935 ;
        RECT 72.380 -10.160 72.700 -10.115 ;
        RECT 73.050 -10.160 73.280 -10.035 ;
        RECT 65.910 -10.405 66.640 -10.235 ;
        RECT 65.910 -10.475 66.140 -10.405 ;
        RECT 57.400 -11.545 59.030 -11.105 ;
        RECT 56.070 -11.965 56.330 -11.925 ;
        RECT 57.710 -11.965 58.710 -11.545 ;
        RECT 62.480 -11.965 62.800 -11.955 ;
        RECT 56.070 -12.205 62.800 -11.965 ;
        RECT 56.070 -12.245 56.330 -12.205 ;
        RECT 57.710 -12.355 58.710 -12.205 ;
        RECT 62.480 -12.215 62.800 -12.205 ;
        RECT 63.050 -13.175 63.320 -10.755 ;
        RECT 64.080 -10.855 65.935 -10.635 ;
        RECT 65.645 -10.865 65.935 -10.855 ;
        RECT 66.445 -11.055 66.615 -10.405 ;
        RECT 70.400 -10.735 71.400 -10.185 ;
        RECT 71.690 -10.615 71.910 -10.185 ;
        RECT 72.380 -10.330 73.280 -10.160 ;
        RECT 72.380 -10.375 72.700 -10.330 ;
        RECT 72.960 -10.360 73.280 -10.330 ;
        RECT 73.050 -10.455 73.280 -10.360 ;
        RECT 73.520 -10.215 73.750 -10.035 ;
        RECT 73.520 -10.385 74.250 -10.215 ;
        RECT 78.400 -10.225 79.920 -10.005 ;
        RECT 86.210 -9.985 87.210 -9.755 ;
        RECT 87.510 -9.915 89.370 -9.695 ;
        RECT 96.655 -9.715 96.945 -9.685 ;
        RECT 87.510 -9.985 87.730 -9.915 ;
        RECT 80.380 -10.200 80.700 -10.155 ;
        RECT 81.050 -10.200 81.280 -10.075 ;
        RECT 73.520 -10.455 73.750 -10.385 ;
        RECT 64.990 -11.495 66.620 -11.055 ;
        RECT 63.670 -11.965 63.930 -11.925 ;
        RECT 65.300 -11.965 66.300 -11.495 ;
        RECT 70.090 -11.965 70.410 -11.955 ;
        RECT 63.670 -12.205 70.410 -11.965 ;
        RECT 63.670 -12.245 63.930 -12.205 ;
        RECT 65.300 -12.305 66.300 -12.205 ;
        RECT 70.090 -12.215 70.410 -12.205 ;
        RECT 70.730 -13.175 71.000 -10.735 ;
        RECT 71.690 -10.835 73.545 -10.615 ;
        RECT 73.255 -10.845 73.545 -10.835 ;
        RECT 74.055 -11.035 74.225 -10.385 ;
        RECT 78.400 -10.775 79.400 -10.225 ;
        RECT 79.690 -10.655 79.910 -10.225 ;
        RECT 80.380 -10.370 81.280 -10.200 ;
        RECT 80.380 -10.415 80.700 -10.370 ;
        RECT 80.960 -10.400 81.280 -10.370 ;
        RECT 81.050 -10.495 81.280 -10.400 ;
        RECT 81.520 -10.255 81.750 -10.075 ;
        RECT 86.210 -10.205 87.730 -9.985 ;
        RECT 93.800 -10.005 94.800 -9.775 ;
        RECT 95.100 -9.935 96.960 -9.715 ;
        RECT 104.045 -9.745 104.335 -9.715 ;
        RECT 95.100 -10.005 95.320 -9.935 ;
        RECT 88.190 -10.180 88.510 -10.135 ;
        RECT 88.860 -10.180 89.090 -10.055 ;
        RECT 81.520 -10.425 82.250 -10.255 ;
        RECT 81.520 -10.495 81.750 -10.425 ;
        RECT 72.600 -11.475 74.230 -11.035 ;
        RECT 71.470 -11.965 71.730 -11.925 ;
        RECT 72.910 -11.965 73.910 -11.475 ;
        RECT 77.970 -11.965 78.290 -11.955 ;
        RECT 71.470 -12.205 78.290 -11.965 ;
        RECT 71.470 -12.245 71.730 -12.205 ;
        RECT 72.910 -12.285 73.910 -12.205 ;
        RECT 77.970 -12.215 78.290 -12.205 ;
        RECT 78.610 -13.175 78.880 -10.775 ;
        RECT 79.690 -10.875 81.545 -10.655 ;
        RECT 81.255 -10.885 81.545 -10.875 ;
        RECT 82.055 -11.075 82.225 -10.425 ;
        RECT 86.210 -10.755 87.210 -10.205 ;
        RECT 87.500 -10.635 87.720 -10.205 ;
        RECT 88.190 -10.350 89.090 -10.180 ;
        RECT 88.190 -10.395 88.510 -10.350 ;
        RECT 88.770 -10.380 89.090 -10.350 ;
        RECT 88.860 -10.475 89.090 -10.380 ;
        RECT 89.330 -10.235 89.560 -10.055 ;
        RECT 93.800 -10.225 95.320 -10.005 ;
        RECT 101.190 -10.035 102.190 -9.805 ;
        RECT 102.490 -9.965 104.350 -9.745 ;
        RECT 102.490 -10.035 102.710 -9.965 ;
        RECT 95.780 -10.200 96.100 -10.155 ;
        RECT 96.450 -10.200 96.680 -10.075 ;
        RECT 89.330 -10.405 90.060 -10.235 ;
        RECT 89.330 -10.475 89.560 -10.405 ;
        RECT 80.600 -11.515 82.230 -11.075 ;
        RECT 79.450 -11.965 79.710 -11.925 ;
        RECT 80.910 -11.965 81.910 -11.515 ;
        RECT 85.840 -11.965 86.160 -11.955 ;
        RECT 79.450 -12.205 86.160 -11.965 ;
        RECT 79.450 -12.245 79.710 -12.205 ;
        RECT 80.910 -12.325 81.910 -12.205 ;
        RECT 85.840 -12.215 86.160 -12.205 ;
        RECT 86.560 -13.175 86.830 -10.755 ;
        RECT 87.500 -10.855 89.355 -10.635 ;
        RECT 89.065 -10.865 89.355 -10.855 ;
        RECT 89.865 -11.055 90.035 -10.405 ;
        RECT 93.800 -10.775 94.800 -10.225 ;
        RECT 95.090 -10.655 95.310 -10.225 ;
        RECT 95.780 -10.370 96.680 -10.200 ;
        RECT 95.780 -10.415 96.100 -10.370 ;
        RECT 96.360 -10.400 96.680 -10.370 ;
        RECT 96.450 -10.495 96.680 -10.400 ;
        RECT 96.920 -10.255 97.150 -10.075 ;
        RECT 101.190 -10.255 102.710 -10.035 ;
        RECT 103.170 -10.230 103.490 -10.185 ;
        RECT 103.840 -10.230 104.070 -10.105 ;
        RECT 96.920 -10.425 97.650 -10.255 ;
        RECT 96.920 -10.495 97.150 -10.425 ;
        RECT 88.410 -11.495 90.040 -11.055 ;
        RECT 87.110 -11.965 87.370 -11.925 ;
        RECT 88.720 -11.965 89.720 -11.495 ;
        RECT 93.780 -11.965 94.100 -11.955 ;
        RECT 87.110 -12.205 94.100 -11.965 ;
        RECT 87.110 -12.245 87.370 -12.205 ;
        RECT 88.720 -12.305 89.720 -12.205 ;
        RECT 93.780 -12.215 94.100 -12.205 ;
        RECT 94.280 -13.175 94.550 -10.775 ;
        RECT 95.090 -10.875 96.945 -10.655 ;
        RECT 96.655 -10.885 96.945 -10.875 ;
        RECT 97.455 -11.075 97.625 -10.425 ;
        RECT 101.190 -10.805 102.190 -10.255 ;
        RECT 102.480 -10.685 102.700 -10.255 ;
        RECT 103.170 -10.400 104.070 -10.230 ;
        RECT 103.170 -10.445 103.490 -10.400 ;
        RECT 103.750 -10.430 104.070 -10.400 ;
        RECT 103.840 -10.525 104.070 -10.430 ;
        RECT 104.310 -10.285 104.540 -10.105 ;
        RECT 104.310 -10.455 105.040 -10.285 ;
        RECT 104.310 -10.525 104.540 -10.455 ;
        RECT 96.000 -11.515 97.630 -11.075 ;
        RECT 94.980 -11.965 95.240 -11.925 ;
        RECT 96.310 -11.965 97.310 -11.515 ;
        RECT 101.030 -11.965 101.350 -11.955 ;
        RECT 94.980 -12.205 101.350 -11.965 ;
        RECT 94.980 -12.245 95.240 -12.205 ;
        RECT 96.310 -12.325 97.310 -12.205 ;
        RECT 101.030 -12.215 101.350 -12.205 ;
        RECT 101.700 -13.175 101.970 -10.805 ;
        RECT 102.480 -10.905 104.335 -10.685 ;
        RECT 104.045 -10.915 104.335 -10.905 ;
        RECT 104.845 -11.105 105.015 -10.455 ;
        RECT 103.390 -11.545 105.020 -11.105 ;
        RECT 102.250 -11.965 102.510 -11.925 ;
        RECT 103.700 -11.965 104.700 -11.545 ;
        RECT 106.650 -11.965 106.970 -11.955 ;
        RECT 102.250 -12.205 106.970 -11.965 ;
        RECT 102.250 -12.245 102.510 -12.205 ;
        RECT 103.700 -12.355 104.700 -12.205 ;
        RECT 106.650 -12.215 106.970 -12.205 ;
        RECT 53.755 -13.445 101.970 -13.175 ;
        RECT 55.450 -13.475 55.720 -13.445 ;
        RECT 86.560 -13.455 86.830 -13.445 ;
        RECT 94.280 -13.455 94.550 -13.445 ;
        RECT 107.325 -13.930 107.595 -6.225 ;
        RECT 108.130 -7.225 108.300 -6.225 ;
        RECT 109.510 -6.190 109.830 -6.155 ;
        RECT 111.815 -6.190 112.005 -5.685 ;
        RECT 112.470 -5.935 113.470 -5.685 ;
        RECT 109.510 -6.380 112.005 -6.190 ;
        RECT 109.510 -6.415 109.830 -6.380 ;
        RECT 110.495 -6.855 110.785 -6.835 ;
        RECT 108.680 -6.865 110.820 -6.855 ;
        RECT 108.650 -7.045 110.820 -6.865 ;
        RECT 108.650 -7.225 108.860 -7.045 ;
        RECT 110.495 -7.065 110.785 -7.045 ;
        RECT 108.130 -7.405 108.860 -7.225 ;
        RECT 108.140 -7.425 108.860 -7.405 ;
        RECT 108.650 -7.835 108.860 -7.425 ;
        RECT 109.540 -7.390 109.800 -7.325 ;
        RECT 110.290 -7.390 110.520 -7.225 ;
        RECT 109.540 -7.580 110.520 -7.390 ;
        RECT 109.540 -7.645 109.800 -7.580 ;
        RECT 110.290 -7.645 110.520 -7.580 ;
        RECT 110.760 -7.395 110.990 -7.225 ;
        RECT 110.760 -7.565 111.840 -7.395 ;
        RECT 110.760 -7.645 110.990 -7.565 ;
        RECT 110.495 -7.835 110.785 -7.805 ;
        RECT 108.650 -8.025 110.800 -7.835 ;
        RECT 110.495 -8.035 110.785 -8.025 ;
        RECT 109.710 -8.700 111.490 -8.345 ;
        RECT 111.655 -8.700 111.825 -7.565 ;
        RECT 109.710 -8.870 111.825 -8.700 ;
        RECT 109.710 -9.165 111.490 -8.870 ;
        RECT 110.160 -9.915 111.160 -9.165 ;
        RECT 108.770 -11.965 109.030 -11.925 ;
        RECT 110.620 -11.965 110.860 -9.915 ;
        RECT 108.770 -12.205 110.870 -11.965 ;
        RECT 108.770 -12.245 109.030 -12.205 ;
        RECT 52.625 -14.200 107.595 -13.930 ;
        RECT 40.950 -15.310 43.940 -14.290 ;
        RECT 9.940 -16.360 40.600 -16.330 ;
        RECT 40.950 -16.360 41.390 -15.310 ;
        RECT 9.940 -16.770 41.390 -16.360 ;
        RECT 38.430 -16.800 41.390 -16.770 ;
        RECT 114.380 -17.905 114.710 4.110 ;
        RECT 115.330 3.860 116.330 4.110 ;
        RECT 119.245 3.465 121.875 3.725 ;
        RECT 119.245 3.255 119.505 3.465 ;
        RECT 115.045 2.985 119.505 3.255 ;
        RECT 116.715 -14.960 116.985 2.985 ;
        RECT 117.415 -8.340 117.685 2.985 ;
        RECT 119.245 1.415 119.505 2.985 ;
        RECT 122.145 2.945 122.445 4.365 ;
        RECT 123.480 2.975 123.700 8.615 ;
        RECT 135.905 8.790 142.415 9.040 ;
        RECT 125.105 6.955 126.105 7.755 ;
        RECT 124.945 6.635 126.785 6.955 ;
        RECT 124.665 6.175 126.785 6.635 ;
        RECT 132.605 6.385 133.605 7.265 ;
        RECT 124.665 5.235 124.945 6.175 ;
        RECT 132.365 6.045 133.915 6.385 ;
        RECT 125.710 5.915 127.800 5.985 ;
        RECT 125.695 5.705 127.800 5.915 ;
        RECT 125.695 5.685 125.985 5.705 ;
        RECT 125.505 5.235 125.735 5.525 ;
        RECT 124.665 4.955 125.775 5.235 ;
        RECT 125.945 5.170 126.175 5.525 ;
        RECT 126.725 5.170 126.985 5.205 ;
        RECT 125.505 4.525 125.735 4.955 ;
        RECT 125.945 4.920 126.985 5.170 ;
        RECT 125.945 4.525 126.175 4.920 ;
        RECT 126.725 4.885 126.985 4.920 ;
        RECT 125.695 4.325 125.985 4.365 ;
        RECT 127.520 4.325 127.800 5.705 ;
        RECT 132.215 5.805 134.045 6.045 ;
        RECT 132.215 5.585 132.455 5.805 ;
        RECT 133.805 5.655 134.045 5.805 ;
        RECT 132.175 5.325 132.495 5.585 ;
        RECT 133.785 5.395 134.045 5.655 ;
        RECT 125.670 4.045 127.800 4.325 ;
        RECT 126.695 3.480 127.015 3.485 ;
        RECT 124.460 3.230 127.015 3.480 ;
        RECT 124.460 2.975 124.710 3.230 ;
        RECT 126.695 3.225 127.015 3.230 ;
        RECT 122.935 2.945 124.710 2.975 ;
        RECT 122.135 2.865 124.710 2.945 ;
        RECT 120.625 2.745 124.710 2.865 ;
        RECT 120.625 2.675 123.185 2.745 ;
        RECT 120.625 2.565 122.445 2.675 ;
        RECT 120.515 1.415 120.745 2.390 ;
        RECT 119.245 1.155 120.745 1.415 ;
        RECT 120.515 -0.110 120.745 1.155 ;
        RECT 120.955 0.535 121.185 2.390 ;
        RECT 122.135 1.055 122.435 2.565 ;
        RECT 124.460 1.115 124.710 2.745 ;
        RECT 127.520 2.695 127.800 4.045 ;
        RECT 131.175 4.945 133.235 5.125 ;
        RECT 131.175 2.825 131.355 4.945 ;
        RECT 132.215 4.675 132.455 4.705 ;
        RECT 132.205 4.355 132.465 4.675 ;
        RECT 133.055 4.545 133.235 4.945 ;
        RECT 132.215 4.065 132.465 4.355 ;
        RECT 132.625 4.315 133.625 4.545 ;
        RECT 132.215 4.055 132.455 4.065 ;
        RECT 132.625 3.875 133.625 4.105 ;
        RECT 133.785 4.035 134.035 5.395 ;
        RECT 134.295 4.755 134.885 5.105 ;
        RECT 133.335 3.130 133.515 3.875 ;
        RECT 134.295 3.755 135.625 4.755 ;
        RECT 134.295 3.305 134.885 3.755 ;
        RECT 135.905 3.130 136.155 8.790 ;
        RECT 138.520 7.465 139.520 8.285 ;
        RECT 138.240 7.195 140.130 7.465 ;
        RECT 138.155 6.865 140.130 7.195 ;
        RECT 138.155 5.775 138.395 6.865 ;
        RECT 138.950 6.325 141.260 6.625 ;
        RECT 138.835 5.775 139.065 6.165 ;
        RECT 138.155 5.535 139.065 5.775 ;
        RECT 138.835 5.165 139.065 5.535 ;
        RECT 139.275 5.700 139.505 6.165 ;
        RECT 139.760 5.700 140.080 5.725 ;
        RECT 139.275 5.490 140.080 5.700 ;
        RECT 139.275 5.165 139.505 5.490 ;
        RECT 139.760 5.465 140.080 5.490 ;
        RECT 140.960 5.015 141.260 6.325 ;
        RECT 138.940 4.715 141.260 5.015 ;
        RECT 139.760 4.020 140.080 4.045 ;
        RECT 137.685 3.810 140.080 4.020 ;
        RECT 137.685 3.685 137.895 3.810 ;
        RECT 139.760 3.785 140.080 3.810 ;
        RECT 133.305 2.880 136.155 3.130 ;
        RECT 137.000 3.425 137.895 3.685 ;
        RECT 129.395 2.695 131.355 2.825 ;
        RECT 127.450 2.665 131.355 2.695 ;
        RECT 125.650 2.645 131.355 2.665 ;
        RECT 125.650 2.465 129.585 2.645 ;
        RECT 125.650 2.385 127.800 2.465 ;
        RECT 125.725 2.365 126.015 2.385 ;
        RECT 125.535 1.115 125.765 2.160 ;
        RECT 122.135 0.755 123.165 1.055 ;
        RECT 124.455 0.865 125.765 1.115 ;
        RECT 120.955 0.275 122.545 0.535 ;
        RECT 120.955 -0.110 121.185 0.275 ;
        RECT 120.705 -0.385 120.995 -0.315 ;
        RECT 122.865 -0.385 123.165 0.755 ;
        RECT 125.535 -0.340 125.765 0.865 ;
        RECT 125.975 0.600 126.205 2.160 ;
        RECT 127.520 0.805 127.800 2.385 ;
        RECT 127.130 0.600 127.390 0.665 ;
        RECT 125.975 0.410 127.390 0.600 ;
        RECT 125.975 -0.340 126.205 0.410 ;
        RECT 127.130 0.345 127.390 0.410 ;
        RECT 127.560 0.175 127.800 0.805 ;
        RECT 120.645 -0.685 123.165 -0.385 ;
        RECT 127.520 -0.495 127.800 0.175 ;
        RECT 125.720 -0.775 127.800 -0.495 ;
        RECT 119.905 -1.415 121.745 -0.825 ;
        RECT 119.905 -1.675 122.545 -1.415 ;
        RECT 124.995 -1.515 126.815 -1.045 ;
        RECT 127.100 -1.515 127.420 -1.480 ;
        RECT 119.905 -1.685 121.745 -1.675 ;
        RECT 120.385 -3.075 121.385 -1.685 ;
        RECT 124.995 -1.705 127.420 -1.515 ;
        RECT 124.995 -1.735 126.815 -1.705 ;
        RECT 125.455 -3.295 126.455 -1.735 ;
        RECT 127.100 -1.740 127.420 -1.705 ;
        RECT 123.215 -3.945 123.565 -3.305 ;
        RECT 122.375 -4.225 124.245 -3.945 ;
        RECT 121.355 -4.775 123.385 -4.555 ;
        RECT 121.355 -6.685 121.575 -4.775 ;
        RECT 122.405 -5.555 122.685 -4.945 ;
        RECT 123.165 -5.055 123.385 -4.775 ;
        RECT 122.835 -5.285 123.835 -5.055 ;
        RECT 124.000 -5.245 124.205 -4.225 ;
        RECT 124.445 -4.935 124.855 -4.515 ;
        RECT 122.835 -5.725 123.835 -5.495 ;
        RECT 123.995 -5.535 124.225 -5.245 ;
        RECT 124.000 -5.585 124.205 -5.535 ;
        RECT 118.965 -6.905 121.575 -6.685 ;
        RECT 123.225 -6.755 123.425 -5.725 ;
        RECT 124.445 -5.935 125.785 -4.935 ;
        RECT 124.445 -6.275 124.855 -5.935 ;
        RECT 128.380 -6.755 128.580 2.465 ;
        RECT 129.395 0.275 129.575 2.465 ;
        RECT 130.315 1.865 131.175 2.295 ;
        RECT 129.735 0.865 131.175 1.865 ;
        RECT 133.335 1.785 133.515 2.880 ;
        RECT 131.445 1.035 131.745 1.595 ;
        RECT 131.920 1.555 134.420 1.785 ;
        RECT 131.920 1.115 134.420 1.345 ;
        RECT 130.315 0.585 131.175 0.865 ;
        RECT 131.985 0.275 132.165 1.115 ;
        RECT 129.395 0.095 132.165 0.275 ;
        RECT 134.565 -0.235 134.865 1.625 ;
        RECT 131.415 -0.535 134.865 -0.235 ;
        RECT 133.155 -1.175 133.465 -0.535 ;
        RECT 118.965 -8.340 119.185 -6.905 ;
        RECT 123.225 -6.955 128.580 -6.755 ;
        RECT 120.365 -7.805 121.165 -7.525 ;
        RECT 117.415 -8.610 119.185 -8.340 ;
        RECT 118.965 -9.435 119.185 -8.610 ;
        RECT 119.505 -8.805 121.165 -7.805 ;
        RECT 123.225 -7.925 123.425 -6.955 ;
        RECT 121.525 -8.765 121.815 -8.085 ;
        RECT 121.960 -8.155 124.460 -7.925 ;
        RECT 124.700 -8.115 124.990 -8.070 ;
        RECT 121.960 -8.595 124.460 -8.365 ;
        RECT 124.665 -8.405 124.990 -8.115 ;
        RECT 120.365 -9.225 121.165 -8.805 ;
        RECT 122.345 -9.435 122.565 -8.595 ;
        RECT 118.965 -9.655 122.565 -9.435 ;
        RECT 124.700 -10.190 124.990 -8.405 ;
        RECT 137.000 -8.835 137.260 3.425 ;
        RECT 137.685 1.735 137.895 3.425 ;
        RECT 140.960 3.465 141.260 4.715 ;
        RECT 142.165 3.695 142.415 8.790 ;
        RECT 158.170 8.235 158.490 10.620 ;
        RECT 144.155 7.125 145.155 7.865 ;
        RECT 157.730 7.245 158.730 8.235 ;
        RECT 143.725 6.665 145.485 7.125 ;
        RECT 157.330 6.985 159.110 7.245 ;
        RECT 143.715 6.465 145.485 6.665 ;
        RECT 143.715 5.375 143.915 6.465 ;
        RECT 152.020 6.280 152.280 6.345 ;
        RECT 152.805 6.280 153.025 6.905 ;
        RECT 157.120 6.665 159.110 6.985 ;
        RECT 144.455 5.935 146.475 6.215 ;
        RECT 152.020 6.090 153.820 6.280 ;
        RECT 152.020 6.025 152.280 6.090 ;
        RECT 144.315 5.375 144.545 5.785 ;
        RECT 143.655 5.175 144.545 5.375 ;
        RECT 144.315 4.785 144.545 5.175 ;
        RECT 144.755 5.285 144.985 5.785 ;
        RECT 145.225 5.285 145.545 5.335 ;
        RECT 144.755 5.125 145.545 5.285 ;
        RECT 144.755 4.785 144.985 5.125 ;
        RECT 145.225 5.075 145.545 5.125 ;
        RECT 144.505 4.615 144.795 4.625 ;
        RECT 146.185 4.615 146.475 5.935 ;
        RECT 150.775 5.495 152.995 5.695 ;
        RECT 150.775 5.245 150.975 5.495 ;
        RECT 150.775 5.155 150.985 5.245 ;
        RECT 144.475 4.575 146.485 4.615 ;
        RECT 144.475 4.335 146.505 4.575 ;
        RECT 145.225 3.825 145.545 3.875 ;
        RECT 142.165 3.515 142.680 3.695 ;
        RECT 143.345 3.665 145.545 3.825 ;
        RECT 143.345 3.515 143.505 3.665 ;
        RECT 145.225 3.615 145.545 3.665 ;
        RECT 146.225 3.695 146.505 4.335 ;
        RECT 150.785 3.895 150.985 5.155 ;
        RECT 152.020 4.915 152.280 5.235 ;
        RECT 152.795 5.125 152.995 5.495 ;
        RECT 152.035 4.645 152.265 4.915 ;
        RECT 152.425 4.895 153.425 5.125 ;
        RECT 153.630 4.935 153.820 6.090 ;
        RECT 152.425 4.455 153.425 4.685 ;
        RECT 153.585 4.645 153.820 4.935 ;
        RECT 153.630 4.620 153.820 4.645 ;
        RECT 154.110 5.195 154.760 5.665 ;
        RECT 157.120 5.625 157.340 6.665 ;
        RECT 158.040 6.155 160.300 6.415 ;
        RECT 157.870 5.625 158.100 5.995 ;
        RECT 157.110 5.405 158.100 5.625 ;
        RECT 147.590 3.695 147.770 3.705 ;
        RECT 148.995 3.695 150.985 3.895 ;
        RECT 142.165 3.465 143.515 3.515 ;
        RECT 140.960 3.275 143.515 3.465 ;
        RECT 146.225 3.455 149.210 3.695 ;
        RECT 152.855 3.685 153.045 4.455 ;
        RECT 154.110 4.195 155.590 5.195 ;
        RECT 157.870 4.995 158.100 5.405 ;
        RECT 158.310 5.620 158.540 5.995 ;
        RECT 158.980 5.620 159.300 5.645 ;
        RECT 158.310 5.410 159.300 5.620 ;
        RECT 158.310 4.995 158.540 5.410 ;
        RECT 158.980 5.385 159.300 5.410 ;
        RECT 158.060 4.825 158.350 4.835 ;
        RECT 160.040 4.825 160.300 6.155 ;
        RECT 157.980 4.565 160.320 4.825 ;
        RECT 154.110 3.895 154.760 4.195 ;
        RECT 158.980 3.890 159.300 3.915 ;
        RECT 155.125 3.685 155.835 3.700 ;
        RECT 140.960 3.215 142.680 3.275 ;
        RECT 140.960 3.185 141.380 3.215 ;
        RECT 140.960 3.005 141.260 3.185 ;
        RECT 139.040 2.705 141.260 3.005 ;
        RECT 138.895 1.735 139.125 2.530 ;
        RECT 137.680 1.525 139.125 1.735 ;
        RECT 138.895 0.030 139.125 1.525 ;
        RECT 139.335 0.535 139.565 2.530 ;
        RECT 140.475 0.555 140.795 0.565 ;
        RECT 140.035 0.535 140.795 0.555 ;
        RECT 139.335 0.315 140.795 0.535 ;
        RECT 139.335 0.295 140.285 0.315 ;
        RECT 140.475 0.305 140.795 0.315 ;
        RECT 139.335 0.030 139.565 0.295 ;
        RECT 140.960 -0.175 141.260 2.705 ;
        RECT 143.345 1.565 143.505 3.275 ;
        RECT 146.225 2.955 146.505 3.455 ;
        RECT 144.485 2.715 146.505 2.955 ;
        RECT 144.345 1.565 144.575 2.520 ;
        RECT 143.345 1.405 144.575 1.565 ;
        RECT 144.345 0.020 144.575 1.405 ;
        RECT 144.785 0.415 145.015 2.520 ;
        RECT 145.685 0.415 146.005 0.440 ;
        RECT 144.785 0.205 146.005 0.415 ;
        RECT 144.785 0.020 145.015 0.205 ;
        RECT 145.685 0.180 146.005 0.205 ;
        RECT 146.225 -0.155 146.505 2.715 ;
        RECT 139.000 -0.475 141.260 -0.175 ;
        RECT 144.535 -0.395 146.505 -0.155 ;
        RECT 144.535 -0.415 144.825 -0.395 ;
        RECT 138.325 -1.135 140.055 -0.735 ;
        RECT 143.695 -1.120 145.435 -0.655 ;
        RECT 145.685 -1.120 146.005 -1.095 ;
        RECT 138.325 -1.395 140.325 -1.135 ;
        RECT 143.695 -1.330 146.005 -1.120 ;
        RECT 138.325 -1.595 140.055 -1.395 ;
        RECT 143.695 -1.595 145.435 -1.330 ;
        RECT 145.685 -1.355 146.005 -1.330 ;
        RECT 138.755 -2.825 139.755 -1.595 ;
        RECT 144.155 -2.635 145.155 -1.595 ;
        RECT 142.595 -4.655 142.915 -4.645 ;
        RECT 143.175 -4.655 144.175 -3.325 ;
        RECT 142.595 -4.895 144.455 -4.655 ;
        RECT 142.595 -4.905 142.915 -4.895 ;
        RECT 141.655 -5.615 143.615 -5.415 ;
        RECT 141.655 -7.435 141.855 -5.615 ;
        RECT 143.415 -5.805 143.615 -5.615 ;
        RECT 142.625 -6.335 142.885 -5.835 ;
        RECT 143.025 -6.035 144.025 -5.805 ;
        RECT 144.215 -5.995 144.455 -4.895 ;
        RECT 143.025 -6.475 144.025 -6.245 ;
        RECT 144.185 -6.285 144.455 -5.995 ;
        RECT 144.215 -6.295 144.455 -6.285 ;
        RECT 144.715 -5.695 145.455 -5.355 ;
        RECT 143.535 -7.365 143.715 -6.475 ;
        RECT 144.715 -6.695 146.245 -5.695 ;
        RECT 144.715 -6.945 145.455 -6.695 ;
        RECT 147.590 -7.365 147.770 3.455 ;
        RECT 148.995 0.795 149.195 3.455 ;
        RECT 152.850 3.430 155.835 3.685 ;
        RECT 156.615 3.680 159.300 3.890 ;
        RECT 156.615 3.465 156.825 3.680 ;
        RECT 158.980 3.655 159.300 3.680 ;
        RECT 152.850 3.420 155.300 3.430 ;
        RECT 150.400 2.415 150.920 2.795 ;
        RECT 149.610 1.395 150.920 2.415 ;
        RECT 152.855 2.265 153.045 3.420 ;
        RECT 150.400 1.225 150.920 1.395 ;
        RECT 150.575 0.795 150.835 0.855 ;
        RECT 148.995 0.595 150.835 0.795 ;
        RECT 150.575 0.535 150.835 0.595 ;
        RECT 151.185 0.345 151.445 2.115 ;
        RECT 151.620 2.035 154.120 2.265 ;
        RECT 154.355 2.075 154.615 2.135 ;
        RECT 151.620 1.595 154.120 1.825 ;
        RECT 154.325 1.785 154.615 2.075 ;
        RECT 151.955 1.445 152.155 1.595 ;
        RECT 151.925 1.125 152.185 1.445 ;
        RECT 154.355 0.345 154.615 1.785 ;
        RECT 151.175 0.045 154.655 0.345 ;
        RECT 151.185 0.025 151.445 0.045 ;
        RECT 152.875 -0.575 153.125 0.045 ;
        RECT 152.455 -1.605 153.455 -0.575 ;
        RECT 141.605 -7.585 141.875 -7.435 ;
        RECT 139.715 -7.775 141.875 -7.585 ;
        RECT 143.535 -7.545 147.770 -7.365 ;
        RECT 139.715 -7.785 141.665 -7.775 ;
        RECT 139.715 -8.835 139.915 -7.785 ;
        RECT 140.975 -8.515 141.565 -8.375 ;
        RECT 137.000 -9.095 139.930 -8.835 ;
        RECT 121.495 -10.480 124.990 -10.190 ;
        RECT 139.715 -10.205 139.915 -9.095 ;
        RECT 140.085 -9.515 141.565 -8.515 ;
        RECT 143.535 -8.645 143.715 -7.545 ;
        RECT 155.565 -8.230 155.835 3.430 ;
        RECT 156.045 3.175 156.830 3.465 ;
        RECT 156.615 1.285 156.825 3.175 ;
        RECT 160.060 3.045 160.320 4.565 ;
        RECT 160.630 3.080 161.630 3.315 ;
        RECT 183.450 3.080 183.710 15.750 ;
        RECT 160.630 3.045 183.710 3.080 ;
        RECT 160.040 2.820 183.710 3.045 ;
        RECT 160.040 2.805 161.630 2.820 ;
        RECT 157.990 2.755 161.630 2.805 ;
        RECT 157.990 2.545 160.320 2.755 ;
        RECT 158.040 2.525 158.330 2.545 ;
        RECT 157.850 1.285 158.080 2.320 ;
        RECT 156.570 1.075 158.080 1.285 ;
        RECT 157.850 -0.180 158.080 1.075 ;
        RECT 158.290 0.175 158.520 2.320 ;
        RECT 159.410 0.175 159.730 0.190 ;
        RECT 158.290 -0.055 159.730 0.175 ;
        RECT 158.290 -0.180 158.520 -0.055 ;
        RECT 159.410 -0.070 159.730 -0.055 ;
        RECT 160.060 -0.345 160.320 2.545 ;
        RECT 160.630 2.285 161.630 2.755 ;
        RECT 157.990 -0.605 160.320 -0.345 ;
        RECT 158.040 -0.615 158.330 -0.605 ;
        RECT 157.320 -1.370 159.130 -0.915 ;
        RECT 159.410 -1.370 159.730 -1.355 ;
        RECT 157.320 -1.600 159.730 -1.370 ;
        RECT 157.320 -1.785 159.130 -1.600 ;
        RECT 159.410 -1.615 159.730 -1.600 ;
        RECT 157.730 -3.135 158.730 -1.785 ;
        RECT 157.980 -3.985 158.310 -3.135 ;
        RECT 163.445 -3.985 163.775 1.695 ;
        RECT 157.980 -4.315 163.775 -3.985 ;
        RECT 157.980 -4.350 158.310 -4.315 ;
        RECT 146.515 -8.500 155.835 -8.230 ;
        RECT 141.825 -9.215 142.155 -8.785 ;
        RECT 142.310 -8.875 144.810 -8.645 ;
        RECT 145.045 -8.835 145.245 -8.825 ;
        RECT 141.860 -9.515 142.120 -9.215 ;
        RECT 142.310 -9.315 144.810 -9.085 ;
        RECT 145.015 -9.125 145.245 -8.835 ;
        RECT 140.975 -9.825 141.565 -9.515 ;
        RECT 142.835 -10.205 143.035 -9.315 ;
        RECT 139.715 -10.405 143.035 -10.205 ;
        RECT 123.085 -10.905 123.405 -10.480 ;
        RECT 141.860 -10.755 142.120 -10.695 ;
        RECT 143.485 -10.755 143.795 -10.745 ;
        RECT 145.045 -10.755 145.245 -9.125 ;
        RECT 122.695 -11.935 123.695 -10.905 ;
        RECT 141.860 -10.955 145.245 -10.755 ;
        RECT 141.860 -11.015 142.120 -10.955 ;
        RECT 143.485 -11.385 143.795 -10.955 ;
        RECT 116.715 -15.030 143.660 -14.960 ;
        RECT 146.515 -15.030 146.785 -8.500 ;
        RECT 116.715 -15.230 146.785 -15.030 ;
        RECT 143.285 -15.300 146.785 -15.230 ;
        RECT 5.375 -18.235 114.710 -17.905 ;
      LAYER met2 ;
        RECT 88.090 86.880 88.530 86.910 ;
        RECT 88.090 86.440 90.205 86.880 ;
        RECT 88.090 86.410 88.530 86.440 ;
        RECT 76.010 76.120 76.530 76.150 ;
        RECT 76.010 75.600 80.815 76.120 ;
        RECT 76.010 75.570 76.530 75.600 ;
        RECT 75.430 61.320 76.430 61.350 ;
        RECT 75.430 60.320 81.950 61.320 ;
        RECT 75.430 60.290 76.430 60.320 ;
        RECT 62.535 52.330 63.005 52.350 ;
        RECT 62.510 51.810 65.210 52.330 ;
        RECT 62.535 51.790 63.005 51.810 ;
        RECT 71.750 50.840 72.270 55.210 ;
        RECT 71.720 50.320 72.300 50.840 ;
        RECT 67.400 35.900 67.920 35.930 ;
        RECT 65.475 35.380 67.920 35.900 ;
        RECT 67.400 35.350 67.920 35.380 ;
        RECT 141.455 32.935 141.785 32.965 ;
        RECT 141.455 32.605 163.775 32.935 ;
        RECT 141.455 32.575 141.785 32.605 ;
        RECT 107.730 32.030 108.050 32.290 ;
        RECT 107.790 30.790 107.990 32.030 ;
        RECT 107.730 30.530 108.050 30.790 ;
        RECT 128.065 29.955 128.355 31.815 ;
        RECT 156.665 31.660 156.985 31.920 ;
        RECT 156.725 30.420 156.925 31.660 ;
        RECT 156.665 30.160 156.985 30.420 ;
        RECT 128.035 29.665 128.385 29.955 ;
        RECT 106.965 27.170 107.285 27.430 ;
        RECT 106.995 25.920 107.255 27.170 ;
        RECT 155.900 26.800 156.220 27.060 ;
        RECT 127.165 26.280 127.505 26.560 ;
        RECT 127.195 25.220 127.475 26.280 ;
        RECT 155.930 25.550 156.190 26.800 ;
        RECT 90.180 22.630 90.440 22.950 ;
        RECT 122.490 22.755 122.750 23.075 ;
        RECT 109.585 22.690 109.845 22.730 ;
        RECT 90.195 21.405 90.425 22.630 ;
        RECT 103.905 22.370 104.165 22.690 ;
        RECT 109.125 22.450 109.845 22.690 ;
        RECT 90.180 21.085 90.440 21.405 ;
        RECT 103.930 21.155 104.140 22.370 ;
        RECT 103.905 20.835 104.165 21.155 ;
        RECT 109.125 21.030 109.365 22.450 ;
        RECT 109.585 22.410 109.845 22.450 ;
        RECT 15.190 20.550 15.510 20.810 ;
        RECT 99.015 20.710 99.335 20.740 ;
        RECT 109.115 20.710 109.375 21.030 ;
        RECT 15.220 19.440 15.480 20.550 ;
        RECT 97.725 20.510 99.335 20.710 ;
        RECT 97.725 20.150 97.925 20.510 ;
        RECT 99.015 20.480 99.335 20.510 ;
        RECT 118.135 20.240 118.435 21.870 ;
        RECT 122.525 20.930 122.715 22.755 ;
        RECT 122.460 20.670 122.780 20.930 ;
        RECT 127.365 20.740 127.625 23.010 ;
        RECT 139.115 22.260 139.375 22.580 ;
        RECT 158.520 22.320 158.780 22.360 ;
        RECT 139.130 21.035 139.360 22.260 ;
        RECT 152.840 22.000 153.100 22.320 ;
        RECT 158.060 22.080 158.780 22.320 ;
        RECT 139.115 20.715 139.375 21.035 ;
        RECT 152.865 20.785 153.075 22.000 ;
        RECT 152.840 20.465 153.100 20.785 ;
        RECT 158.060 20.660 158.300 22.080 ;
        RECT 158.520 22.040 158.780 22.080 ;
        RECT 147.950 20.340 148.270 20.370 ;
        RECT 158.050 20.340 158.310 20.660 ;
        RECT 97.665 19.890 97.985 20.150 ;
        RECT 118.105 19.940 118.465 20.240 ;
        RECT 146.660 20.140 148.270 20.340 ;
        RECT 146.660 19.780 146.860 20.140 ;
        RECT 147.950 20.110 148.270 20.140 ;
        RECT 16.490 19.730 16.750 19.760 ;
        RECT 16.490 19.470 18.060 19.730 ;
        RECT 146.600 19.520 146.920 19.780 ;
        RECT 16.490 19.440 16.750 19.470 ;
        RECT 25.565 18.615 25.895 18.645 ;
        RECT 25.565 18.285 30.005 18.615 ;
        RECT 25.565 18.255 25.895 18.285 ;
        RECT 16.930 17.720 17.190 18.040 ;
        RECT 3.780 16.230 4.040 16.550 ;
        RECT 16.980 16.430 17.140 17.720 ;
        RECT 24.800 16.500 25.060 16.820 ;
        RECT 3.810 15.470 4.010 16.230 ;
        RECT 16.900 16.170 17.220 16.430 ;
        RECT 3.780 15.150 4.040 15.470 ;
        RECT 24.825 15.245 25.035 16.500 ;
        RECT 26.760 16.100 27.080 16.360 ;
        RECT 28.780 16.310 29.100 16.570 ;
        RECT 55.255 16.345 55.585 19.355 ;
        RECT 122.895 17.790 123.155 18.110 ;
        RECT 90.610 17.360 90.870 17.680 ;
        RECT 104.365 17.400 104.625 17.720 ;
        RECT 24.800 14.925 25.060 15.245 ;
        RECT -22.610 14.330 -22.290 14.590 ;
        RECT -22.550 11.920 -22.350 14.330 ;
        RECT -10.330 14.300 -10.070 14.620 ;
        RECT 11.380 14.610 12.890 14.870 ;
        RECT 26.805 14.450 27.035 16.100 ;
        RECT 28.850 15.340 29.030 16.310 ;
        RECT 90.635 15.950 90.845 17.360 ;
        RECT 97.570 16.100 97.890 16.360 ;
        RECT 104.415 16.260 104.575 17.400 ;
        RECT 109.830 17.230 110.090 17.550 ;
        RECT 90.610 15.630 90.870 15.950 ;
        RECT 28.810 15.020 29.070 15.340 ;
        RECT 97.635 15.250 97.825 16.100 ;
        RECT 104.365 15.940 104.625 16.260 ;
        RECT 109.855 15.870 110.065 17.230 ;
        RECT 117.385 16.660 117.705 16.920 ;
        RECT 117.425 16.010 117.665 16.660 ;
        RECT 122.900 16.390 123.150 17.790 ;
        RECT 122.865 16.130 123.185 16.390 ;
        RECT 109.830 15.550 110.090 15.870 ;
        RECT 117.415 15.690 117.675 16.010 ;
        RECT 128.035 15.810 128.295 17.870 ;
        RECT 139.545 16.990 139.805 17.310 ;
        RECT 153.300 17.030 153.560 17.350 ;
        RECT 139.570 15.580 139.780 16.990 ;
        RECT 146.505 15.730 146.825 15.990 ;
        RECT 153.350 15.890 153.510 17.030 ;
        RECT 158.765 16.860 159.025 17.180 ;
        RECT 139.545 15.260 139.805 15.580 ;
        RECT 97.570 14.990 97.890 15.250 ;
        RECT 146.570 14.880 146.760 15.730 ;
        RECT 153.300 15.570 153.560 15.890 ;
        RECT 158.790 15.500 159.000 16.860 ;
        RECT 158.765 15.180 159.025 15.500 ;
        RECT 146.505 14.620 146.825 14.880 ;
        RECT -10.300 12.140 -10.100 14.300 ;
        RECT 26.760 14.190 27.080 14.450 ;
        RECT 14.360 14.010 14.620 14.090 ;
        RECT 15.520 14.010 15.840 14.060 ;
        RECT -1.220 13.680 -0.960 13.740 ;
        RECT 0.000 13.680 0.320 13.710 ;
        RECT -1.220 13.480 0.320 13.680 ;
        RECT 4.240 13.650 4.500 13.970 ;
        RECT 14.360 13.850 15.840 14.010 ;
        RECT 14.360 13.770 14.620 13.850 ;
        RECT 15.520 13.800 15.840 13.850 ;
        RECT -1.220 13.420 -0.960 13.480 ;
        RECT 0.000 13.450 0.320 13.480 ;
        RECT 4.260 12.580 4.480 13.650 ;
        RECT 55.225 13.295 55.615 13.625 ;
        RECT 4.240 12.260 4.500 12.580 ;
        RECT -22.580 11.600 -22.320 11.920 ;
        RECT -10.360 11.880 -10.040 12.140 ;
        RECT -22.590 9.860 -22.310 9.895 ;
        RECT -21.550 9.860 -21.250 11.140 ;
        RECT -10.905 10.385 -10.585 10.645 ;
        RECT 11.930 10.420 12.210 10.450 ;
        RECT -22.600 9.560 -21.250 9.860 ;
        RECT -15.030 9.750 -14.770 10.070 ;
        RECT -22.590 9.525 -22.310 9.560 ;
        RECT -15.000 9.210 -14.800 9.750 ;
        RECT -23.150 9.010 -14.800 9.210 ;
        RECT -23.150 8.290 -22.950 9.010 ;
        RECT -19.700 8.470 -19.500 9.010 ;
        RECT -15.000 8.470 -14.800 9.010 ;
        RECT -22.600 8.290 -22.300 8.355 ;
        RECT -23.210 8.030 -22.890 8.290 ;
        RECT -22.610 8.030 -22.290 8.290 ;
        RECT -19.730 8.150 -19.470 8.470 ;
        RECT -15.030 8.150 -14.770 8.470 ;
        RECT -22.600 7.965 -22.300 8.030 ;
        RECT -10.840 7.515 -10.645 10.385 ;
        RECT 10.780 10.140 12.210 10.420 ;
        RECT 11.930 10.110 12.210 10.140 ;
        RECT 55.255 8.895 55.585 13.295 ;
        RECT 82.800 12.230 83.240 12.260 ;
        RECT 82.800 11.790 88.920 12.230 ;
        RECT 82.800 11.760 83.240 11.790 ;
        RECT -23.320 7.260 -23.000 7.290 ;
        RECT -16.160 7.260 -15.840 7.290 ;
        RECT -23.320 7.060 -15.840 7.260 ;
        RECT -23.320 7.030 -23.000 7.060 ;
        RECT -16.160 7.030 -15.840 7.060 ;
        RECT -23.225 6.105 -22.965 6.425 ;
        RECT -23.185 4.025 -23.000 6.105 ;
        RECT -12.305 4.505 -11.985 4.545 ;
        RECT -10.835 4.505 -10.650 7.515 ;
        RECT 17.970 7.200 18.290 7.460 ;
        RECT 4.680 6.620 4.940 6.670 ;
        RECT 6.150 6.620 6.470 6.640 ;
        RECT 4.680 6.400 6.470 6.620 ;
        RECT 4.680 6.350 4.940 6.400 ;
        RECT 6.150 6.380 6.470 6.400 ;
        RECT 9.020 6.620 9.280 6.670 ;
        RECT 10.810 6.620 11.130 6.640 ;
        RECT 9.020 6.400 11.130 6.620 ;
        RECT 9.020 6.350 9.280 6.400 ;
        RECT 10.810 6.380 11.130 6.400 ;
        RECT 18.030 5.790 18.230 7.200 ;
        RECT 18.000 5.470 18.260 5.790 ;
        RECT -12.305 4.320 -10.650 4.505 ;
        RECT -12.305 4.285 -11.985 4.320 ;
        RECT -23.220 3.705 -22.960 4.025 ;
        RECT -21.030 2.950 -20.770 3.270 ;
        RECT -21.010 0.650 -20.790 2.950 ;
        RECT -14.030 2.800 -13.770 3.120 ;
        RECT -21.710 0.230 -21.390 0.490 ;
        RECT -21.650 -1.030 -21.450 0.230 ;
        RECT -21.680 -1.350 -21.420 -1.030 ;
        RECT -21.000 -1.730 -20.800 0.650 ;
        RECT -20.560 -1.310 -20.240 -1.280 ;
        RECT -19.940 -1.310 -18.000 -1.290 ;
        RECT -20.560 -1.490 -18.000 -1.310 ;
        RECT -20.560 -1.510 -19.790 -1.490 ;
        RECT -20.560 -1.540 -20.240 -1.510 ;
        RECT -29.910 -1.990 -29.590 -1.960 ;
        RECT -28.480 -1.990 -28.220 -1.930 ;
        RECT -29.910 -2.190 -28.220 -1.990 ;
        RECT -21.030 -2.050 -20.770 -1.730 ;
        RECT -29.910 -2.220 -29.590 -2.190 ;
        RECT -28.480 -2.250 -28.220 -2.190 ;
        RECT -24.900 -3.490 -20.950 -3.290 ;
        RECT -24.900 -4.310 -24.700 -3.490 ;
        RECT -21.150 -4.180 -20.950 -3.490 ;
        RECT -18.200 -4.110 -18.000 -1.490 ;
        RECT -24.960 -4.570 -24.640 -4.310 ;
        RECT -21.180 -4.500 -20.920 -4.180 ;
        RECT -18.260 -4.370 -17.940 -4.110 ;
        RECT -14.000 -4.160 -13.800 2.800 ;
        RECT -11.530 2.470 -11.270 2.535 ;
        RECT -10.835 2.470 -10.650 4.320 ;
        RECT 2.355 3.955 2.765 4.305 ;
        RECT -0.640 3.785 -0.290 3.815 ;
        RECT 2.385 3.785 2.735 3.955 ;
        RECT -0.640 3.435 2.735 3.785 ;
        RECT 44.420 3.460 44.760 6.150 ;
        RECT 151.990 6.055 152.310 6.315 ;
        RECT 121.585 3.435 121.845 5.495 ;
        RECT 132.205 5.295 132.465 5.615 ;
        RECT 139.790 5.435 140.050 5.755 ;
        RECT 126.695 4.915 127.015 5.175 ;
        RECT 126.730 3.515 126.980 4.915 ;
        RECT 132.215 4.645 132.455 5.295 ;
        RECT 132.175 4.385 132.495 4.645 ;
        RECT 139.815 4.075 140.025 5.435 ;
        RECT 145.255 5.045 145.515 5.365 ;
        RECT 152.055 5.205 152.245 6.055 ;
        RECT 159.010 5.355 159.270 5.675 ;
        RECT 139.790 3.755 140.050 4.075 ;
        RECT 145.305 3.905 145.465 5.045 ;
        RECT 151.990 4.945 152.310 5.205 ;
        RECT 159.035 3.945 159.245 5.355 ;
        RECT 145.255 3.585 145.515 3.905 ;
        RECT 159.010 3.625 159.270 3.945 ;
        RECT -0.640 3.405 -0.290 3.435 ;
        RECT 126.725 3.195 126.985 3.515 ;
        RECT -11.530 2.285 -10.650 2.470 ;
        RECT 4.820 2.400 5.080 2.720 ;
        RECT 35.930 2.450 36.190 2.770 ;
        RECT -11.530 2.215 -11.270 2.285 ;
        RECT -10.835 0.705 -10.650 2.285 ;
        RECT 4.850 1.620 5.050 2.400 ;
        RECT 4.820 1.300 5.080 1.620 ;
        RECT 35.955 1.480 36.165 2.450 ;
        RECT 107.100 1.740 107.500 2.080 ;
        RECT 35.930 1.160 36.190 1.480 ;
        RECT 12.070 0.810 13.600 1.090 ;
        RECT -10.835 0.520 -9.910 0.705 ;
        RECT -10.090 -1.030 -9.920 0.520 ;
        RECT -9.230 0.250 -8.970 0.570 ;
        RECT 20.170 0.440 20.490 0.700 ;
        RECT 107.130 0.540 107.470 1.740 ;
        RECT 163.445 1.665 163.775 32.605 ;
        RECT 177.000 29.585 177.290 31.445 ;
        RECT 176.970 29.295 177.320 29.585 ;
        RECT 176.100 25.910 176.440 26.190 ;
        RECT 176.130 24.850 176.410 25.910 ;
        RECT 171.425 22.385 171.685 22.705 ;
        RECT 167.070 19.870 167.370 21.500 ;
        RECT 171.460 20.560 171.650 22.385 ;
        RECT 171.395 20.300 171.715 20.560 ;
        RECT 176.300 20.370 176.560 22.640 ;
        RECT 167.040 19.570 167.400 19.870 ;
        RECT 171.830 17.420 172.090 17.740 ;
        RECT 166.320 16.290 166.640 16.550 ;
        RECT 166.360 15.640 166.600 16.290 ;
        RECT 171.835 16.020 172.085 17.420 ;
        RECT 171.800 15.760 172.120 16.020 ;
        RECT 166.350 15.320 166.610 15.640 ;
        RECT 176.970 15.440 177.230 17.500 ;
        RECT 131.415 1.065 131.775 1.365 ;
        RECT 151.895 1.155 152.215 1.415 ;
        RECT 163.415 1.335 163.805 1.665 ;
        RECT -9.200 -1.010 -9.000 0.250 ;
        RECT 15.440 0.230 15.700 0.300 ;
        RECT 16.360 0.230 16.680 0.270 ;
        RECT 15.440 0.050 16.680 0.230 ;
        RECT 15.440 -0.020 15.700 0.050 ;
        RECT 16.360 0.010 16.680 0.050 ;
        RECT 20.240 -0.330 20.420 0.440 ;
        RECT 53.430 0.310 53.690 0.355 ;
        RECT 55.800 0.310 56.120 0.325 ;
        RECT 53.430 0.080 56.120 0.310 ;
        RECT 53.430 0.035 53.690 0.080 ;
        RECT 55.800 0.065 56.120 0.080 ;
        RECT 61.990 0.310 62.250 0.355 ;
        RECT 63.490 0.310 63.810 0.325 ;
        RECT 61.990 0.080 63.810 0.310 ;
        RECT 61.990 0.035 62.250 0.080 ;
        RECT 63.490 0.065 63.810 0.080 ;
        RECT 69.810 0.310 70.070 0.355 ;
        RECT 70.930 0.310 71.250 0.325 ;
        RECT 69.810 0.080 71.250 0.310 ;
        RECT 69.810 0.035 70.070 0.080 ;
        RECT 70.930 0.065 71.250 0.080 ;
        RECT 77.730 0.310 78.050 0.325 ;
        RECT 78.850 0.310 79.170 0.325 ;
        RECT 77.730 0.080 79.170 0.310 ;
        RECT 77.730 0.065 78.050 0.080 ;
        RECT 78.850 0.065 79.170 0.080 ;
        RECT 85.400 0.310 85.660 0.355 ;
        RECT 86.720 0.310 87.040 0.325 ;
        RECT 85.400 0.080 87.040 0.310 ;
        RECT 85.400 0.035 85.660 0.080 ;
        RECT 86.720 0.065 87.040 0.080 ;
        RECT 93.330 0.310 93.590 0.355 ;
        RECT 94.480 0.310 94.800 0.325 ;
        RECT 93.330 0.080 94.800 0.310 ;
        RECT 93.330 0.035 93.590 0.080 ;
        RECT 94.480 0.065 94.800 0.080 ;
        RECT 100.560 0.310 100.820 0.355 ;
        RECT 101.580 0.310 101.900 0.325 ;
        RECT 100.560 0.080 101.900 0.310 ;
        RECT 100.560 0.035 100.820 0.080 ;
        RECT 101.580 0.065 101.900 0.080 ;
        RECT 20.200 -0.650 20.460 -0.330 ;
        RECT 4.980 -0.940 5.300 -0.680 ;
        RECT 56.810 -0.735 57.070 -0.415 ;
        RECT 64.400 -0.685 64.660 -0.365 ;
        RECT 72.010 -0.665 72.270 -0.345 ;
        RECT -10.135 -1.350 -9.875 -1.030 ;
        RECT -9.260 -1.270 -8.940 -1.010 ;
        RECT 5.045 -1.710 5.235 -0.940 ;
        RECT 15.310 -1.190 15.630 -0.930 ;
        RECT 0.500 -2.040 0.760 -1.980 ;
        RECT 1.800 -2.040 2.120 -2.010 ;
        RECT 5.010 -2.030 5.270 -1.710 ;
        RECT 15.380 -1.870 15.560 -1.190 ;
        RECT 0.500 -2.240 2.120 -2.040 ;
        RECT 15.340 -2.190 15.600 -1.870 ;
        RECT 56.820 -1.955 57.060 -0.735 ;
        RECT 56.820 -2.205 57.370 -1.955 ;
        RECT 58.760 -2.050 59.020 -1.730 ;
        RECT 64.410 -1.905 64.650 -0.685 ;
        RECT 57.050 -2.215 57.370 -2.205 ;
        RECT 0.500 -2.300 0.760 -2.240 ;
        RECT 1.800 -2.270 2.120 -2.240 ;
        RECT -13.030 -2.900 -12.770 -2.580 ;
        RECT -14.060 -4.420 -13.740 -4.160 ;
        RECT -13.000 -4.260 -12.800 -2.900 ;
        RECT 58.805 -3.265 58.975 -2.050 ;
        RECT 64.410 -2.155 64.960 -1.905 ;
        RECT 66.350 -2.000 66.610 -1.680 ;
        RECT 72.020 -1.885 72.260 -0.665 ;
        RECT 80.010 -0.705 80.270 -0.385 ;
        RECT 87.820 -0.685 88.080 -0.365 ;
        RECT 64.640 -2.165 64.960 -2.155 ;
        RECT 66.395 -3.215 66.565 -2.000 ;
        RECT 72.020 -2.135 72.570 -1.885 ;
        RECT 73.960 -1.980 74.220 -1.660 ;
        RECT 80.020 -1.925 80.260 -0.705 ;
        RECT 72.250 -2.145 72.570 -2.135 ;
        RECT 74.005 -3.195 74.175 -1.980 ;
        RECT 80.020 -2.175 80.570 -1.925 ;
        RECT 81.960 -2.020 82.220 -1.700 ;
        RECT 87.830 -1.905 88.070 -0.685 ;
        RECT 95.410 -0.705 95.670 -0.385 ;
        RECT 80.250 -2.185 80.570 -2.175 ;
        RECT 57.460 -3.405 58.975 -3.265 ;
        RECT 12.130 -4.180 12.450 -4.175 ;
        RECT 13.240 -4.180 13.500 -4.145 ;
        RECT -13.060 -4.520 -12.740 -4.260 ;
        RECT 12.130 -4.430 13.500 -4.180 ;
        RECT 12.130 -4.435 12.450 -4.430 ;
        RECT 13.240 -4.465 13.500 -4.430 ;
        RECT 57.460 -4.755 57.600 -3.405 ;
        RECT 58.805 -3.420 58.975 -3.405 ;
        RECT 65.050 -3.355 66.565 -3.215 ;
        RECT 65.050 -4.705 65.190 -3.355 ;
        RECT 66.395 -3.370 66.565 -3.355 ;
        RECT 72.660 -3.335 74.175 -3.195 ;
        RECT 82.005 -3.235 82.175 -2.020 ;
        RECT 87.830 -2.155 88.380 -1.905 ;
        RECT 89.770 -2.000 90.030 -1.680 ;
        RECT 95.420 -1.925 95.660 -0.705 ;
        RECT 102.800 -0.735 103.060 -0.415 ;
        RECT 88.060 -2.165 88.380 -2.155 ;
        RECT 89.815 -3.215 89.985 -2.000 ;
        RECT 95.420 -2.175 95.970 -1.925 ;
        RECT 97.360 -2.020 97.620 -1.700 ;
        RECT 102.810 -1.955 103.050 -0.735 ;
        RECT 122.255 -1.705 122.515 0.565 ;
        RECT 127.100 0.375 127.420 0.635 ;
        RECT 127.165 -1.450 127.355 0.375 ;
        RECT 131.445 -0.565 131.745 1.065 ;
        RECT 150.545 0.795 150.865 0.825 ;
        RECT 151.955 0.795 152.155 1.155 ;
        RECT 150.545 0.595 152.155 0.795 ;
        RECT 140.505 0.275 140.765 0.595 ;
        RECT 150.545 0.565 150.865 0.595 ;
        RECT 140.035 -1.145 140.295 -1.105 ;
        RECT 140.515 -1.145 140.755 0.275 ;
        RECT 145.715 0.150 145.975 0.470 ;
        RECT 145.740 -1.065 145.950 0.150 ;
        RECT 159.440 -0.100 159.700 0.220 ;
        RECT 140.035 -1.385 140.755 -1.145 ;
        RECT 145.715 -1.385 145.975 -1.065 ;
        RECT 159.455 -1.325 159.685 -0.100 ;
        RECT 140.035 -1.425 140.295 -1.385 ;
        RECT 95.650 -2.185 95.970 -2.175 ;
        RECT 72.660 -4.685 72.800 -3.335 ;
        RECT 74.005 -3.350 74.175 -3.335 ;
        RECT 80.660 -3.375 82.175 -3.235 ;
        RECT 57.400 -5.075 57.660 -4.755 ;
        RECT 64.990 -5.025 65.250 -4.705 ;
        RECT 72.600 -5.005 72.860 -4.685 ;
        RECT 80.660 -4.725 80.800 -3.375 ;
        RECT 82.005 -3.390 82.175 -3.375 ;
        RECT 88.470 -3.355 89.985 -3.215 ;
        RECT 97.405 -3.235 97.575 -2.020 ;
        RECT 102.810 -2.205 103.360 -1.955 ;
        RECT 104.750 -2.050 105.010 -1.730 ;
        RECT 127.130 -1.770 127.390 -1.450 ;
        RECT 159.440 -1.645 159.700 -1.325 ;
        RECT 103.040 -2.215 103.360 -2.205 ;
        RECT 88.470 -4.705 88.610 -3.355 ;
        RECT 89.815 -3.370 89.985 -3.355 ;
        RECT 96.060 -3.375 97.575 -3.235 ;
        RECT 104.795 -3.265 104.965 -2.050 ;
        RECT 109.340 -2.895 109.600 -2.575 ;
        RECT 80.600 -5.045 80.860 -4.725 ;
        RECT 88.410 -5.025 88.670 -4.705 ;
        RECT 96.060 -4.725 96.200 -3.375 ;
        RECT 97.405 -3.390 97.575 -3.375 ;
        RECT 103.450 -3.405 104.965 -3.265 ;
        RECT 96.000 -5.045 96.260 -4.725 ;
        RECT 103.450 -4.755 103.590 -3.405 ;
        RECT 104.795 -3.420 104.965 -3.405 ;
        RECT 109.380 -4.085 109.560 -2.895 ;
        RECT 109.310 -4.345 109.630 -4.085 ;
        RECT 103.390 -5.075 103.650 -4.755 ;
        RECT 122.405 -4.975 122.685 -3.915 ;
        RECT 122.375 -5.255 122.715 -4.975 ;
        RECT 142.625 -5.865 142.885 -4.615 ;
        RECT 142.595 -6.125 142.915 -5.865 ;
        RECT 20.200 -6.490 20.460 -6.170 ;
        RECT 109.540 -6.445 109.800 -6.125 ;
        RECT 5.430 -6.840 5.710 -6.810 ;
        RECT 10.000 -6.840 10.275 -6.810 ;
        RECT 5.430 -7.115 7.115 -6.840 ;
        RECT 10.000 -7.115 11.395 -6.840 ;
        RECT 5.430 -7.150 5.710 -7.115 ;
        RECT 10.000 -7.145 10.275 -7.115 ;
        RECT 20.240 -7.450 20.420 -6.490 ;
        RECT 57.110 -7.005 57.370 -6.685 ;
        RECT 64.700 -6.955 64.960 -6.635 ;
        RECT 72.310 -6.935 72.570 -6.615 ;
        RECT 20.200 -7.770 20.460 -7.450 ;
        RECT 48.450 -7.455 48.710 -7.135 ;
        RECT 48.475 -8.345 48.685 -7.455 ;
        RECT 57.150 -7.705 57.330 -7.005 ;
        RECT 64.740 -7.655 64.920 -6.955 ;
        RECT 72.350 -7.635 72.530 -6.935 ;
        RECT 80.310 -6.975 80.570 -6.655 ;
        RECT 88.120 -6.955 88.380 -6.635 ;
        RECT 57.080 -7.965 57.400 -7.705 ;
        RECT 64.670 -7.915 64.990 -7.655 ;
        RECT 72.280 -7.895 72.600 -7.635 ;
        RECT 80.350 -7.675 80.530 -6.975 ;
        RECT 88.160 -7.655 88.340 -6.955 ;
        RECT 95.710 -6.975 95.970 -6.655 ;
        RECT 80.280 -7.935 80.600 -7.675 ;
        RECT 88.090 -7.915 88.410 -7.655 ;
        RECT 95.750 -7.675 95.930 -6.975 ;
        RECT 103.100 -7.005 103.360 -6.685 ;
        RECT 95.680 -7.935 96.000 -7.675 ;
        RECT 103.140 -7.705 103.320 -7.005 ;
        RECT 109.575 -7.355 109.765 -6.445 ;
        RECT 109.510 -7.615 109.830 -7.355 ;
        RECT 103.070 -7.965 103.390 -7.705 ;
        RECT 48.450 -8.665 48.710 -8.345 ;
        RECT 121.495 -8.650 121.845 -8.360 ;
        RECT 29.085 -9.420 29.405 -9.160 ;
        RECT 29.150 -10.330 29.340 -9.420 ;
        RECT 57.210 -9.635 57.470 -9.315 ;
        RECT 64.800 -9.585 65.060 -9.265 ;
        RECT 72.410 -9.565 72.670 -9.245 ;
        RECT 57.255 -10.155 57.425 -9.635 ;
        RECT 64.845 -10.105 65.015 -9.585 ;
        RECT 72.455 -10.085 72.625 -9.565 ;
        RECT 80.410 -9.605 80.670 -9.285 ;
        RECT 88.220 -9.585 88.480 -9.265 ;
        RECT 29.115 -10.650 29.375 -10.330 ;
        RECT 57.210 -10.475 57.470 -10.155 ;
        RECT 64.800 -10.425 65.060 -10.105 ;
        RECT 72.410 -10.405 72.670 -10.085 ;
        RECT 80.455 -10.125 80.625 -9.605 ;
        RECT 88.265 -10.105 88.435 -9.585 ;
        RECT 95.810 -9.605 96.070 -9.285 ;
        RECT 80.410 -10.445 80.670 -10.125 ;
        RECT 88.220 -10.425 88.480 -10.105 ;
        RECT 95.855 -10.125 96.025 -9.605 ;
        RECT 103.200 -9.635 103.460 -9.315 ;
        RECT 95.810 -10.445 96.070 -10.125 ;
        RECT 103.245 -10.155 103.415 -9.635 ;
        RECT 103.200 -10.475 103.460 -10.155 ;
        RECT 121.525 -10.510 121.815 -8.650 ;
        RECT 141.830 -9.485 142.150 -9.225 ;
        RECT 46.470 -10.600 46.810 -10.570 ;
        RECT 46.470 -10.940 48.450 -10.600 ;
        RECT 141.890 -10.725 142.090 -9.485 ;
        RECT 46.470 -10.970 46.810 -10.940 ;
        RECT 141.830 -10.985 142.150 -10.725 ;
        RECT 52.080 -11.965 52.340 -11.925 ;
        RECT 53.270 -11.965 53.590 -11.955 ;
        RECT 52.080 -12.205 53.590 -11.965 ;
        RECT 52.080 -12.245 52.340 -12.205 ;
        RECT 53.270 -12.215 53.590 -12.205 ;
        RECT 54.940 -11.965 55.200 -11.925 ;
        RECT 56.040 -11.965 56.360 -11.955 ;
        RECT 54.940 -12.205 56.360 -11.965 ;
        RECT 54.940 -12.245 55.200 -12.205 ;
        RECT 56.040 -12.215 56.360 -12.205 ;
        RECT 62.510 -11.965 62.770 -11.925 ;
        RECT 63.640 -11.965 63.960 -11.955 ;
        RECT 62.510 -12.205 63.960 -11.965 ;
        RECT 62.510 -12.245 62.770 -12.205 ;
        RECT 63.640 -12.215 63.960 -12.205 ;
        RECT 70.120 -11.965 70.380 -11.925 ;
        RECT 71.440 -11.965 71.760 -11.955 ;
        RECT 70.120 -12.205 71.760 -11.965 ;
        RECT 70.120 -12.245 70.380 -12.205 ;
        RECT 71.440 -12.215 71.760 -12.205 ;
        RECT 78.000 -11.965 78.260 -11.925 ;
        RECT 79.420 -11.965 79.740 -11.955 ;
        RECT 78.000 -12.205 79.740 -11.965 ;
        RECT 78.000 -12.245 78.260 -12.205 ;
        RECT 79.420 -12.215 79.740 -12.205 ;
        RECT 85.870 -11.965 86.130 -11.925 ;
        RECT 87.080 -11.965 87.400 -11.955 ;
        RECT 85.870 -12.205 87.400 -11.965 ;
        RECT 85.870 -12.245 86.130 -12.205 ;
        RECT 87.080 -12.215 87.400 -12.205 ;
        RECT 93.810 -11.965 94.070 -11.925 ;
        RECT 94.950 -11.965 95.270 -11.955 ;
        RECT 93.810 -12.205 95.270 -11.965 ;
        RECT 93.810 -12.245 94.070 -12.205 ;
        RECT 94.950 -12.215 95.270 -12.205 ;
        RECT 101.060 -11.965 101.320 -11.925 ;
        RECT 102.220 -11.965 102.540 -11.955 ;
        RECT 101.060 -12.205 102.540 -11.965 ;
        RECT 101.060 -12.245 101.320 -12.205 ;
        RECT 102.220 -12.215 102.540 -12.205 ;
        RECT 106.680 -11.965 106.940 -11.925 ;
        RECT 108.740 -11.965 109.060 -11.955 ;
        RECT 106.680 -12.205 109.060 -11.965 ;
        RECT 106.680 -12.245 106.940 -12.205 ;
        RECT 108.740 -12.215 109.060 -12.205 ;
        RECT 53.785 -13.175 54.055 -13.145 ;
        RECT 51.095 -13.445 54.055 -13.175 ;
        RECT 53.785 -13.475 54.055 -13.445 ;
      LAYER met3 ;
        RECT -319.110 399.070 -288.710 430.930 ;
        RECT -287.510 399.070 -257.110 430.930 ;
        RECT -255.910 399.070 -225.510 430.930 ;
        RECT -224.310 399.070 -193.910 430.930 ;
        RECT -192.710 399.070 -162.310 430.930 ;
        RECT -161.110 399.070 -130.710 430.930 ;
        RECT -129.510 399.070 -99.110 430.930 ;
        RECT -97.910 399.070 -67.510 430.930 ;
        RECT -66.310 399.070 -35.910 430.930 ;
        RECT -34.710 399.070 -4.310 430.930 ;
        RECT -3.110 399.070 27.290 430.930 ;
        RECT 28.490 399.070 58.890 430.930 ;
        RECT -321.670 381.205 -321.150 384.170 ;
        RECT -321.695 380.695 -321.125 381.205 ;
        RECT -321.670 380.690 -321.150 380.695 ;
        RECT -319.110 366.010 -288.710 397.870 ;
        RECT -287.510 366.010 -257.110 397.870 ;
        RECT -255.910 366.010 -225.510 397.870 ;
        RECT -224.310 366.010 -193.910 397.870 ;
        RECT -192.710 366.010 -162.310 397.870 ;
        RECT -161.110 366.010 -130.710 397.870 ;
        RECT -129.510 366.010 -99.110 397.870 ;
        RECT -97.910 366.010 -67.510 397.870 ;
        RECT -66.310 366.010 -35.910 397.870 ;
        RECT -34.710 366.010 -4.310 397.870 ;
        RECT -3.110 366.010 27.290 397.870 ;
        RECT 28.490 366.010 58.890 397.870 ;
        RECT -319.110 332.950 -288.710 364.810 ;
        RECT -287.510 332.950 -257.110 364.810 ;
        RECT -255.910 332.950 -225.510 364.810 ;
        RECT -224.310 332.950 -193.910 364.810 ;
        RECT -192.710 332.950 -162.310 364.810 ;
        RECT -161.110 332.950 -130.710 364.810 ;
        RECT -129.510 332.950 -99.110 364.810 ;
        RECT -97.910 332.950 -67.510 364.810 ;
        RECT -66.310 332.950 -35.910 364.810 ;
        RECT -34.710 332.950 -4.310 364.810 ;
        RECT -3.110 332.950 27.290 364.810 ;
        RECT 28.490 332.950 58.890 364.810 ;
        RECT 59.910 347.630 60.430 351.200 ;
        RECT 59.915 347.605 60.425 347.630 ;
        RECT -320.800 315.425 -320.280 317.700 ;
        RECT -320.825 314.915 -320.255 315.425 ;
        RECT -320.800 314.910 -320.280 314.915 ;
        RECT -319.110 299.890 -288.710 331.750 ;
        RECT -287.510 299.890 -257.110 331.750 ;
        RECT -255.910 299.890 -225.510 331.750 ;
        RECT -224.310 299.890 -193.910 331.750 ;
        RECT -192.710 299.890 -162.310 331.750 ;
        RECT -161.110 299.890 -130.710 331.750 ;
        RECT -129.510 299.890 -99.110 331.750 ;
        RECT -97.910 299.890 -67.510 331.750 ;
        RECT -66.310 299.890 -35.910 331.750 ;
        RECT -34.710 299.890 -4.310 331.750 ;
        RECT -3.110 299.890 27.290 331.750 ;
        RECT 28.490 299.890 58.890 331.750 ;
        RECT -319.110 266.830 -288.710 298.690 ;
        RECT -287.510 266.830 -257.110 298.690 ;
        RECT -255.910 266.830 -225.510 298.690 ;
        RECT -224.310 266.830 -193.910 298.690 ;
        RECT -192.710 266.830 -162.310 298.690 ;
        RECT -161.110 266.830 -130.710 298.690 ;
        RECT -129.510 266.830 -99.110 298.690 ;
        RECT -97.910 266.830 -67.510 298.690 ;
        RECT -66.310 266.830 -35.910 298.690 ;
        RECT -34.710 266.830 -4.310 298.690 ;
        RECT -3.110 266.830 27.290 298.690 ;
        RECT 28.490 266.830 58.890 298.690 ;
        RECT 59.960 282.345 60.480 285.680 ;
        RECT 59.935 281.835 60.505 282.345 ;
        RECT 59.960 281.830 60.480 281.835 ;
        RECT -320.950 249.295 -320.430 251.720 ;
        RECT -320.975 248.785 -320.405 249.295 ;
        RECT -320.950 248.780 -320.430 248.785 ;
        RECT -319.110 233.770 -288.710 265.630 ;
        RECT -287.510 233.770 -257.110 265.630 ;
        RECT -255.910 233.770 -225.510 265.630 ;
        RECT -224.310 233.770 -193.910 265.630 ;
        RECT -192.710 233.770 -162.310 265.630 ;
        RECT -161.110 233.770 -130.710 265.630 ;
        RECT -129.510 233.770 -99.110 265.630 ;
        RECT -97.910 233.770 -67.510 265.630 ;
        RECT -66.310 233.770 -35.910 265.630 ;
        RECT -34.710 233.770 -4.310 265.630 ;
        RECT -3.110 233.770 27.290 265.630 ;
        RECT 28.490 233.770 58.890 265.630 ;
        RECT -319.110 200.710 -288.710 232.570 ;
        RECT -287.510 200.710 -257.110 232.570 ;
        RECT -255.910 200.710 -225.510 232.570 ;
        RECT -224.310 200.710 -193.910 232.570 ;
        RECT -192.710 200.710 -162.310 232.570 ;
        RECT -161.110 200.710 -130.710 232.570 ;
        RECT -129.510 200.710 -99.110 232.570 ;
        RECT -97.910 200.710 -67.510 232.570 ;
        RECT -66.310 200.710 -35.910 232.570 ;
        RECT -34.710 200.710 -4.310 232.570 ;
        RECT -3.110 200.710 27.290 232.570 ;
        RECT 28.490 200.710 58.890 232.570 ;
        RECT 60.000 216.105 60.520 218.870 ;
        RECT 59.975 215.595 60.545 216.105 ;
        RECT 60.000 215.590 60.520 215.595 ;
        RECT 95.865 202.740 99.735 202.745 ;
        RECT 95.840 202.215 99.735 202.740 ;
        RECT 100.940 202.220 131.340 234.080 ;
        RECT 132.540 202.220 162.940 234.080 ;
        RECT 164.140 202.220 194.540 234.080 ;
        RECT 195.740 202.220 226.140 234.080 ;
        RECT 227.340 202.220 257.740 234.080 ;
        RECT 95.865 202.210 99.735 202.215 ;
        RECT -321.350 182.710 -320.830 185.800 ;
        RECT -321.345 182.685 -320.835 182.710 ;
        RECT -319.110 167.650 -288.710 199.510 ;
        RECT -287.510 167.650 -257.110 199.510 ;
        RECT -255.910 167.650 -225.510 199.510 ;
        RECT -224.310 167.650 -193.910 199.510 ;
        RECT -192.710 167.650 -162.310 199.510 ;
        RECT -161.110 167.650 -130.710 199.510 ;
        RECT -129.510 167.650 -99.110 199.510 ;
        RECT -97.910 167.650 -67.510 199.510 ;
        RECT -66.310 167.650 -35.910 199.510 ;
        RECT -34.710 167.650 -4.310 199.510 ;
        RECT -3.110 167.650 27.290 199.510 ;
        RECT 28.490 167.650 58.890 199.510 ;
        RECT 100.940 169.160 131.340 201.020 ;
        RECT 132.540 169.160 162.940 201.020 ;
        RECT 164.140 169.160 194.540 201.020 ;
        RECT 195.740 169.160 226.140 201.020 ;
        RECT 227.340 169.160 257.740 201.020 ;
        RECT 259.100 171.420 259.680 171.940 ;
        RECT -319.110 134.590 -288.710 166.450 ;
        RECT -287.510 134.590 -257.110 166.450 ;
        RECT -255.910 134.590 -225.510 166.450 ;
        RECT -224.310 134.590 -193.910 166.450 ;
        RECT -192.710 134.590 -162.310 166.450 ;
        RECT -161.110 134.590 -130.710 166.450 ;
        RECT -129.510 134.590 -99.110 166.450 ;
        RECT -97.910 134.590 -67.510 166.450 ;
        RECT -66.310 134.590 -35.910 166.450 ;
        RECT -34.710 134.590 -4.310 166.450 ;
        RECT -3.110 134.590 27.290 166.450 ;
        RECT 28.490 134.590 58.890 166.450 ;
        RECT 60.190 150.185 60.710 152.760 ;
        RECT 60.165 149.675 60.735 150.185 ;
        RECT 60.190 149.670 60.710 149.675 ;
        RECT 100.940 136.100 131.340 167.960 ;
        RECT 132.540 136.100 162.940 167.960 ;
        RECT 164.140 136.100 194.540 167.960 ;
        RECT 195.740 136.100 226.140 167.960 ;
        RECT 227.340 136.100 257.740 167.960 ;
        RECT 259.130 167.615 259.650 171.420 ;
        RECT 259.105 167.105 259.675 167.615 ;
        RECT 259.130 167.100 259.650 167.105 ;
        RECT -321.130 117.155 -320.610 119.670 ;
        RECT -321.155 116.645 -320.585 117.155 ;
        RECT -321.130 116.640 -320.610 116.645 ;
        RECT -319.110 101.530 -288.710 133.390 ;
        RECT -287.510 101.530 -257.110 133.390 ;
        RECT -255.910 101.530 -225.510 133.390 ;
        RECT -224.310 101.530 -193.910 133.390 ;
        RECT -192.710 101.530 -162.310 133.390 ;
        RECT -161.110 101.530 -130.710 133.390 ;
        RECT -129.510 101.530 -99.110 133.390 ;
        RECT -97.910 101.530 -67.510 133.390 ;
        RECT -66.310 101.530 -35.910 133.390 ;
        RECT -34.710 101.530 -4.310 133.390 ;
        RECT -3.110 101.530 27.290 133.390 ;
        RECT 28.490 101.530 58.890 133.390 ;
        RECT 98.750 118.395 99.270 121.500 ;
        RECT 98.725 117.885 99.295 118.395 ;
        RECT 98.750 117.880 99.270 117.885 ;
        RECT 100.940 103.040 131.340 134.900 ;
        RECT 132.540 103.040 162.940 134.900 ;
        RECT 164.140 103.040 194.540 134.900 ;
        RECT 195.740 103.040 226.140 134.900 ;
        RECT 227.340 103.040 257.740 134.900 ;
        RECT 258.710 103.575 261.920 103.580 ;
        RECT 258.710 103.065 261.945 103.575 ;
        RECT 258.710 103.060 261.920 103.065 ;
        RECT -319.110 68.470 -288.710 100.330 ;
        RECT -287.510 68.470 -257.110 100.330 ;
        RECT -255.910 68.470 -225.510 100.330 ;
        RECT -224.310 68.470 -193.910 100.330 ;
        RECT -192.710 68.470 -162.310 100.330 ;
        RECT -161.110 68.470 -130.710 100.330 ;
        RECT -129.510 68.470 -99.110 100.330 ;
        RECT -97.910 68.470 -67.510 100.330 ;
        RECT -66.310 68.470 -35.910 100.330 ;
        RECT -34.710 68.470 -4.310 100.330 ;
        RECT -3.110 68.470 27.290 100.330 ;
        RECT 28.490 68.470 58.890 100.330 ;
        RECT 89.695 86.880 90.185 86.905 ;
        RECT 60.230 84.115 60.750 86.470 ;
        RECT 89.695 86.440 92.000 86.880 ;
        RECT 89.695 86.415 90.185 86.440 ;
        RECT 60.205 83.605 60.775 84.115 ;
        RECT 60.230 83.600 60.750 83.605 ;
        RECT 80.225 76.120 80.795 76.145 ;
        RECT 80.225 75.600 86.580 76.120 ;
        RECT 80.225 75.575 80.795 75.600 ;
        RECT 100.940 69.980 131.340 101.840 ;
        RECT 132.540 69.980 162.940 101.840 ;
        RECT 164.140 69.980 194.540 101.840 ;
        RECT 195.740 69.980 226.140 101.840 ;
        RECT 227.340 69.980 257.740 101.840 ;
        RECT -322.000 50.815 -321.480 54.420 ;
        RECT -322.025 50.305 -321.455 50.815 ;
        RECT -322.000 50.300 -321.480 50.305 ;
        RECT -319.110 35.410 -288.710 67.270 ;
        RECT -287.510 35.410 -257.110 67.270 ;
        RECT -255.910 35.410 -225.510 67.270 ;
        RECT -224.310 35.410 -193.910 67.270 ;
        RECT -192.710 35.410 -162.310 67.270 ;
        RECT -161.110 35.410 -130.710 67.270 ;
        RECT -129.510 35.410 -99.110 67.270 ;
        RECT -97.910 35.410 -67.510 67.270 ;
        RECT -66.310 35.410 -35.910 67.270 ;
        RECT -34.710 35.410 -4.310 67.270 ;
        RECT -3.110 35.410 27.290 67.270 ;
        RECT 28.490 35.410 58.890 67.270 ;
        RECT 60.255 52.330 60.765 52.355 ;
        RECT 60.250 51.810 63.030 52.330 ;
        RECT 60.255 51.785 60.765 51.810 ;
        RECT 65.495 35.900 66.065 35.925 ;
        RECT 63.000 35.380 66.065 35.900 ;
        RECT 65.495 35.355 66.065 35.380 ;
        RECT -22.615 9.545 -22.285 9.875 ;
        RECT -22.600 8.335 -22.300 9.545 ;
        RECT -22.625 7.985 -22.275 8.335 ;
      LAYER met4 ;
        RECT -324.350 415.990 -319.180 416.050 ;
        RECT -318.715 415.990 -289.105 430.535 ;
        RECT -287.115 415.990 -257.505 430.535 ;
        RECT -255.515 415.990 -225.905 430.535 ;
        RECT -223.915 415.990 -194.305 430.535 ;
        RECT -192.315 415.990 -162.705 430.535 ;
        RECT -160.715 415.990 -131.105 430.535 ;
        RECT -129.115 415.990 -99.505 430.535 ;
        RECT -97.515 415.990 -67.905 430.535 ;
        RECT -65.915 415.990 -36.305 430.535 ;
        RECT -34.315 415.990 -4.705 430.535 ;
        RECT -2.715 415.990 26.895 430.535 ;
        RECT 28.885 415.990 58.495 430.535 ;
        RECT -324.350 415.530 59.490 415.990 ;
        RECT -324.350 382.930 -323.830 415.530 ;
        RECT -319.710 415.470 59.490 415.530 ;
        RECT -318.715 400.925 -289.105 415.470 ;
        RECT -287.115 400.925 -257.505 415.470 ;
        RECT -255.515 400.925 -225.905 415.470 ;
        RECT -223.915 400.925 -194.305 415.470 ;
        RECT -192.315 400.925 -162.705 415.470 ;
        RECT -160.715 400.925 -131.105 415.470 ;
        RECT -129.115 400.925 -99.505 415.470 ;
        RECT -97.515 400.925 -67.905 415.470 ;
        RECT -65.915 400.925 -36.305 415.470 ;
        RECT -34.315 400.925 -4.705 415.470 ;
        RECT -2.715 400.925 26.895 415.470 ;
        RECT 28.885 400.925 58.495 415.470 ;
        RECT -319.710 399.530 59.490 399.590 ;
        RECT -321.670 399.070 59.490 399.530 ;
        RECT -321.670 399.010 -319.270 399.070 ;
        RECT -321.670 384.145 -321.150 399.010 ;
        RECT -321.675 383.615 -321.145 384.145 ;
        RECT -318.715 382.930 -289.105 397.475 ;
        RECT -287.115 382.930 -257.505 397.475 ;
        RECT -255.515 382.930 -225.905 397.475 ;
        RECT -223.915 382.930 -194.305 397.475 ;
        RECT -192.315 382.930 -162.705 397.475 ;
        RECT -160.715 382.930 -131.105 397.475 ;
        RECT -129.115 382.930 -99.505 397.475 ;
        RECT -97.515 382.930 -67.905 397.475 ;
        RECT -65.915 382.930 -36.305 397.475 ;
        RECT -34.315 382.930 -4.705 397.475 ;
        RECT -2.715 382.930 26.895 397.475 ;
        RECT 28.885 382.930 58.495 397.475 ;
        RECT -324.350 382.910 59.490 382.930 ;
        RECT -324.350 382.410 63.020 382.910 ;
        RECT -321.670 366.530 -321.150 381.210 ;
        RECT -318.715 367.865 -289.105 382.410 ;
        RECT -287.115 367.865 -257.505 382.410 ;
        RECT -255.515 367.865 -225.905 382.410 ;
        RECT -223.915 367.865 -194.305 382.410 ;
        RECT -192.315 367.865 -162.705 382.410 ;
        RECT -160.715 367.865 -131.105 382.410 ;
        RECT -129.115 367.865 -99.505 382.410 ;
        RECT -97.515 367.865 -67.905 382.410 ;
        RECT -65.915 367.865 -36.305 382.410 ;
        RECT -34.315 367.865 -4.705 382.410 ;
        RECT -2.715 367.865 26.895 382.410 ;
        RECT 28.885 367.865 58.495 382.410 ;
        RECT 59.030 382.390 63.020 382.410 ;
        RECT -321.670 366.505 59.490 366.530 ;
        RECT -321.670 366.010 60.435 366.505 ;
        RECT 59.025 365.975 60.435 366.010 ;
        RECT -318.715 349.870 -289.105 364.415 ;
        RECT -287.115 349.870 -257.505 364.415 ;
        RECT -255.515 349.870 -225.905 364.415 ;
        RECT -223.915 349.870 -194.305 364.415 ;
        RECT -192.315 349.870 -162.705 364.415 ;
        RECT -160.715 349.870 -131.105 364.415 ;
        RECT -129.115 349.870 -99.505 364.415 ;
        RECT -97.515 349.870 -67.905 364.415 ;
        RECT -65.915 349.870 -36.305 364.415 ;
        RECT -34.315 349.870 -4.705 364.415 ;
        RECT -2.715 349.870 26.895 364.415 ;
        RECT 28.885 349.870 58.495 364.415 ;
        RECT 59.905 350.645 60.435 365.975 ;
        RECT 62.500 349.870 63.020 382.390 ;
        RECT -319.710 349.820 63.020 349.870 ;
        RECT -322.910 349.350 63.020 349.820 ;
        RECT -322.910 349.300 -319.140 349.350 ;
        RECT -322.910 316.810 -322.390 349.300 ;
        RECT -318.715 334.805 -289.105 349.350 ;
        RECT -287.115 334.805 -257.505 349.350 ;
        RECT -255.515 334.805 -225.905 349.350 ;
        RECT -223.915 334.805 -194.305 349.350 ;
        RECT -192.315 334.805 -162.705 349.350 ;
        RECT -160.715 334.805 -131.105 349.350 ;
        RECT -129.115 334.805 -99.505 349.350 ;
        RECT -97.515 334.805 -67.905 349.350 ;
        RECT -65.915 334.805 -36.305 349.350 ;
        RECT -34.315 334.805 -4.705 349.350 ;
        RECT -2.715 334.805 26.895 349.350 ;
        RECT 28.885 334.805 58.495 349.350 ;
        RECT 59.910 333.470 60.430 348.150 ;
        RECT -319.710 333.430 60.430 333.470 ;
        RECT -320.800 332.950 60.430 333.430 ;
        RECT -320.800 332.910 -319.120 332.950 ;
        RECT -320.800 317.675 -320.280 332.910 ;
        RECT -320.805 317.145 -320.275 317.675 ;
        RECT -318.715 316.810 -289.105 331.355 ;
        RECT -287.115 316.810 -257.505 331.355 ;
        RECT -255.515 316.810 -225.905 331.355 ;
        RECT -223.915 316.810 -194.305 331.355 ;
        RECT -192.315 316.810 -162.705 331.355 ;
        RECT -160.715 316.810 -131.105 331.355 ;
        RECT -129.115 316.810 -99.505 331.355 ;
        RECT -97.515 316.810 -67.905 331.355 ;
        RECT -65.915 316.810 -36.305 331.355 ;
        RECT -34.315 316.810 -4.705 331.355 ;
        RECT -2.715 316.810 26.895 331.355 ;
        RECT 28.885 316.810 58.495 331.355 ;
        RECT -322.910 316.770 59.490 316.810 ;
        RECT -322.910 316.290 64.330 316.770 ;
        RECT -320.800 300.410 -320.280 315.430 ;
        RECT -318.715 301.745 -289.105 316.290 ;
        RECT -287.115 301.745 -257.505 316.290 ;
        RECT -255.515 301.745 -225.905 316.290 ;
        RECT -223.915 301.745 -194.305 316.290 ;
        RECT -192.315 301.745 -162.705 316.290 ;
        RECT -160.715 301.745 -131.105 316.290 ;
        RECT -129.115 301.745 -99.505 316.290 ;
        RECT -97.515 301.745 -67.905 316.290 ;
        RECT -65.915 301.745 -36.305 316.290 ;
        RECT -34.315 301.745 -4.705 316.290 ;
        RECT -2.715 301.745 26.895 316.290 ;
        RECT 28.885 301.745 58.495 316.290 ;
        RECT 59.140 316.250 64.330 316.290 ;
        RECT 58.920 300.410 60.480 300.460 ;
        RECT -320.800 299.940 60.480 300.410 ;
        RECT -320.800 299.890 59.490 299.940 ;
        RECT -322.180 283.750 -319.140 283.840 ;
        RECT -318.715 283.750 -289.105 298.295 ;
        RECT -287.115 283.750 -257.505 298.295 ;
        RECT -255.515 283.750 -225.905 298.295 ;
        RECT -223.915 283.750 -194.305 298.295 ;
        RECT -192.315 283.750 -162.705 298.295 ;
        RECT -160.715 283.750 -131.105 298.295 ;
        RECT -129.115 283.750 -99.505 298.295 ;
        RECT -97.515 283.750 -67.905 298.295 ;
        RECT -65.915 283.750 -36.305 298.295 ;
        RECT -34.315 283.750 -4.705 298.295 ;
        RECT -2.715 283.750 26.895 298.295 ;
        RECT 28.885 283.750 58.495 298.295 ;
        RECT 59.960 285.655 60.480 299.940 ;
        RECT 59.955 285.125 60.485 285.655 ;
        RECT 63.810 283.750 64.330 316.250 ;
        RECT -322.180 283.320 64.330 283.750 ;
        RECT -322.180 250.690 -321.660 283.320 ;
        RECT -319.710 283.230 64.330 283.320 ;
        RECT -318.715 268.685 -289.105 283.230 ;
        RECT -287.115 268.685 -257.505 283.230 ;
        RECT -255.515 268.685 -225.905 283.230 ;
        RECT -223.915 268.685 -194.305 283.230 ;
        RECT -192.315 268.685 -162.705 283.230 ;
        RECT -160.715 268.685 -131.105 283.230 ;
        RECT -129.115 268.685 -99.505 283.230 ;
        RECT -97.515 268.685 -67.905 283.230 ;
        RECT -65.915 268.685 -36.305 283.230 ;
        RECT -34.315 268.685 -4.705 283.230 ;
        RECT -2.715 268.685 26.895 283.230 ;
        RECT 28.885 268.685 58.495 283.230 ;
        RECT 59.960 267.350 60.480 282.350 ;
        RECT -319.710 267.250 60.480 267.350 ;
        RECT -320.950 266.830 60.480 267.250 ;
        RECT -320.950 266.730 -319.300 266.830 ;
        RECT -320.950 251.695 -320.430 266.730 ;
        RECT -320.955 251.165 -320.425 251.695 ;
        RECT -318.715 250.690 -289.105 265.235 ;
        RECT -287.115 250.690 -257.505 265.235 ;
        RECT -255.515 250.690 -225.905 265.235 ;
        RECT -223.915 250.690 -194.305 265.235 ;
        RECT -192.315 250.690 -162.705 265.235 ;
        RECT -160.715 250.690 -131.105 265.235 ;
        RECT -129.115 250.690 -99.505 265.235 ;
        RECT -97.515 250.690 -67.905 265.235 ;
        RECT -65.915 250.690 -36.305 265.235 ;
        RECT -34.315 250.690 -4.705 265.235 ;
        RECT -2.715 250.690 26.895 265.235 ;
        RECT 28.885 250.690 58.495 265.235 ;
        RECT 58.980 250.690 63.590 250.730 ;
        RECT -322.180 250.210 63.590 250.690 ;
        RECT -322.180 250.170 59.490 250.210 ;
        RECT -320.950 234.290 -320.430 249.300 ;
        RECT -318.715 235.625 -289.105 250.170 ;
        RECT -287.115 235.625 -257.505 250.170 ;
        RECT -255.515 235.625 -225.905 250.170 ;
        RECT -223.915 235.625 -194.305 250.170 ;
        RECT -192.315 235.625 -162.705 250.170 ;
        RECT -160.715 235.625 -131.105 250.170 ;
        RECT -129.115 235.625 -99.505 250.170 ;
        RECT -97.515 235.625 -67.905 250.170 ;
        RECT -65.915 235.625 -36.305 250.170 ;
        RECT -34.315 235.625 -4.705 250.170 ;
        RECT -2.715 235.625 26.895 250.170 ;
        RECT 28.885 235.625 58.495 250.170 ;
        RECT 59.150 234.290 60.520 234.330 ;
        RECT -320.950 233.810 60.520 234.290 ;
        RECT -320.950 233.770 59.490 233.810 ;
        RECT -318.715 217.630 -289.105 232.175 ;
        RECT -287.115 217.630 -257.505 232.175 ;
        RECT -255.515 217.630 -225.905 232.175 ;
        RECT -223.915 217.630 -194.305 232.175 ;
        RECT -192.315 217.630 -162.705 232.175 ;
        RECT -160.715 217.630 -131.105 232.175 ;
        RECT -129.115 217.630 -99.505 232.175 ;
        RECT -97.515 217.630 -67.905 232.175 ;
        RECT -65.915 217.630 -36.305 232.175 ;
        RECT -34.315 217.630 -4.705 232.175 ;
        RECT -2.715 217.630 26.895 232.175 ;
        RECT 28.885 217.630 58.495 232.175 ;
        RECT 60.000 218.845 60.520 233.810 ;
        RECT 59.995 218.315 60.525 218.845 ;
        RECT 63.070 217.630 63.590 250.210 ;
        RECT 101.335 219.140 130.945 233.685 ;
        RECT 132.935 219.140 162.545 233.685 ;
        RECT 164.535 219.140 194.145 233.685 ;
        RECT 196.135 219.140 225.745 233.685 ;
        RECT 227.735 219.140 257.345 233.685 ;
        RECT 100.340 219.130 258.340 219.140 ;
        RECT -324.520 217.110 63.590 217.630 ;
        RECT 98.210 218.620 258.340 219.130 ;
        RECT 98.210 218.610 130.945 218.620 ;
        RECT -324.520 184.570 -324.000 217.110 ;
        RECT -318.715 202.565 -289.105 217.110 ;
        RECT -287.115 202.565 -257.505 217.110 ;
        RECT -255.515 202.565 -225.905 217.110 ;
        RECT -223.915 202.565 -194.305 217.110 ;
        RECT -192.315 202.565 -162.705 217.110 ;
        RECT -160.715 202.565 -131.105 217.110 ;
        RECT -129.115 202.565 -99.505 217.110 ;
        RECT -97.515 202.565 -67.905 217.110 ;
        RECT -65.915 202.565 -36.305 217.110 ;
        RECT -34.315 202.565 -4.705 217.110 ;
        RECT -2.715 202.565 26.895 217.110 ;
        RECT 28.885 202.565 58.495 217.110 ;
        RECT -321.350 201.230 -318.790 201.260 ;
        RECT 60.000 201.230 60.520 216.110 ;
        RECT -321.350 200.740 60.520 201.230 ;
        RECT -321.350 185.775 -320.830 200.740 ;
        RECT -319.710 200.710 60.520 200.740 ;
        RECT -321.355 185.245 -320.825 185.775 ;
        RECT -318.715 184.570 -289.105 199.115 ;
        RECT -287.115 184.570 -257.505 199.115 ;
        RECT -255.515 184.570 -225.905 199.115 ;
        RECT -223.915 184.570 -194.305 199.115 ;
        RECT -192.315 184.570 -162.705 199.115 ;
        RECT -160.715 184.570 -131.105 199.115 ;
        RECT -129.115 184.570 -99.505 199.115 ;
        RECT -97.515 184.570 -67.905 199.115 ;
        RECT -65.915 184.570 -36.305 199.115 ;
        RECT -34.315 184.570 -4.705 199.115 ;
        RECT -2.715 184.570 26.895 199.115 ;
        RECT 28.885 184.570 58.495 199.115 ;
        RECT 59.020 184.570 62.040 184.580 ;
        RECT -324.520 184.060 62.040 184.570 ;
        RECT -324.520 184.050 59.490 184.060 ;
        RECT -321.350 168.170 -320.830 183.230 ;
        RECT -318.715 169.505 -289.105 184.050 ;
        RECT -287.115 169.505 -257.505 184.050 ;
        RECT -255.515 169.505 -225.905 184.050 ;
        RECT -223.915 169.505 -194.305 184.050 ;
        RECT -192.315 169.505 -162.705 184.050 ;
        RECT -160.715 169.505 -131.105 184.050 ;
        RECT -129.115 169.505 -99.505 184.050 ;
        RECT -97.515 169.505 -67.905 184.050 ;
        RECT -65.915 169.505 -36.305 184.050 ;
        RECT -34.315 169.505 -4.705 184.050 ;
        RECT -2.715 169.505 26.895 184.050 ;
        RECT 28.885 169.505 58.495 184.050 ;
        RECT -321.350 168.110 59.490 168.170 ;
        RECT -321.350 167.650 60.710 168.110 ;
        RECT 59.280 167.590 60.710 167.650 ;
        RECT -318.715 151.510 -289.105 166.055 ;
        RECT -287.115 151.510 -257.505 166.055 ;
        RECT -255.515 151.510 -225.905 166.055 ;
        RECT -223.915 151.510 -194.305 166.055 ;
        RECT -192.315 151.510 -162.705 166.055 ;
        RECT -160.715 151.510 -131.105 166.055 ;
        RECT -129.115 151.510 -99.505 166.055 ;
        RECT -97.515 151.510 -67.905 166.055 ;
        RECT -65.915 151.510 -36.305 166.055 ;
        RECT -34.315 151.510 -4.705 166.055 ;
        RECT -2.715 151.510 26.895 166.055 ;
        RECT 28.885 151.510 58.495 166.055 ;
        RECT 60.190 152.735 60.710 167.590 ;
        RECT 60.185 152.205 60.715 152.735 ;
        RECT 61.520 151.510 62.040 184.060 ;
        RECT 95.865 169.680 96.400 202.745 ;
        RECT 98.210 186.080 98.730 218.610 ;
        RECT 101.335 204.075 130.945 218.610 ;
        RECT 132.935 204.075 162.545 218.620 ;
        RECT 164.535 204.075 194.145 218.620 ;
        RECT 196.135 204.075 225.745 218.620 ;
        RECT 227.735 204.075 257.345 218.620 ;
        RECT 99.165 202.745 99.710 202.750 ;
        RECT 99.165 202.740 100.805 202.745 ;
        RECT 99.165 202.220 258.340 202.740 ;
        RECT 99.165 202.210 100.805 202.220 ;
        RECT 99.165 202.205 99.710 202.210 ;
        RECT 101.335 186.080 130.945 200.625 ;
        RECT 132.935 186.080 162.545 200.625 ;
        RECT 164.535 186.080 194.145 200.625 ;
        RECT 196.135 186.080 225.745 200.625 ;
        RECT 227.735 186.080 257.345 200.625 ;
        RECT 257.930 186.080 259.650 186.100 ;
        RECT 98.210 185.580 259.650 186.080 ;
        RECT 98.210 185.560 258.340 185.580 ;
        RECT 101.335 171.015 130.945 185.560 ;
        RECT 132.935 171.015 162.545 185.560 ;
        RECT 164.535 171.015 194.145 185.560 ;
        RECT 196.135 171.015 225.745 185.560 ;
        RECT 227.735 171.015 257.345 185.560 ;
        RECT 259.130 171.945 259.650 185.580 ;
        RECT 259.125 171.415 259.655 171.945 ;
        RECT 258.045 169.680 261.550 169.685 ;
        RECT 95.865 169.170 261.550 169.680 ;
        RECT 95.865 169.160 258.340 169.170 ;
        RECT 95.865 169.155 96.400 169.160 ;
        RECT 101.335 153.020 130.945 167.565 ;
        RECT 132.935 153.020 162.545 167.565 ;
        RECT 164.535 153.020 194.145 167.565 ;
        RECT 196.135 153.020 225.745 167.565 ;
        RECT 227.735 153.020 257.345 167.565 ;
        RECT 259.130 153.020 259.650 167.620 ;
        RECT 100.340 153.010 259.650 153.020 ;
        RECT -319.710 151.450 62.040 151.510 ;
        RECT -323.040 150.990 62.040 151.450 ;
        RECT 96.610 152.500 259.650 153.010 ;
        RECT 96.610 152.490 100.880 152.500 ;
        RECT -323.040 150.930 -319.160 150.990 ;
        RECT -323.040 118.450 -322.520 150.930 ;
        RECT -318.715 136.445 -289.105 150.990 ;
        RECT -287.115 136.445 -257.505 150.990 ;
        RECT -255.515 136.445 -225.905 150.990 ;
        RECT -223.915 136.445 -194.305 150.990 ;
        RECT -192.315 136.445 -162.705 150.990 ;
        RECT -160.715 136.445 -131.105 150.990 ;
        RECT -129.115 136.445 -99.505 150.990 ;
        RECT -97.515 136.445 -67.905 150.990 ;
        RECT -65.915 136.445 -36.305 150.990 ;
        RECT -34.315 136.445 -4.705 150.990 ;
        RECT -2.715 136.445 26.895 150.990 ;
        RECT 28.885 136.445 58.495 150.990 ;
        RECT -321.130 135.110 -319.290 135.140 ;
        RECT 60.190 135.110 60.710 150.190 ;
        RECT -321.130 134.620 60.710 135.110 ;
        RECT -321.130 119.645 -320.610 134.620 ;
        RECT -319.710 134.590 60.710 134.620 ;
        RECT -321.135 119.115 -320.605 119.645 ;
        RECT -318.715 118.450 -289.105 132.995 ;
        RECT -287.115 118.450 -257.505 132.995 ;
        RECT -255.515 118.450 -225.905 132.995 ;
        RECT -223.915 118.450 -194.305 132.995 ;
        RECT -192.315 118.450 -162.705 132.995 ;
        RECT -160.715 118.450 -131.105 132.995 ;
        RECT -129.115 118.450 -99.505 132.995 ;
        RECT -97.515 118.450 -67.905 132.995 ;
        RECT -65.915 118.450 -36.305 132.995 ;
        RECT -34.315 118.450 -4.705 132.995 ;
        RECT -2.715 118.450 26.895 132.995 ;
        RECT 28.885 118.450 58.495 132.995 ;
        RECT 96.610 119.960 97.130 152.490 ;
        RECT 101.335 137.955 130.945 152.500 ;
        RECT 132.935 137.955 162.545 152.500 ;
        RECT 164.535 137.955 194.145 152.500 ;
        RECT 196.135 137.955 225.745 152.500 ;
        RECT 227.735 137.955 257.345 152.500 ;
        RECT 261.035 136.620 261.550 169.170 ;
        RECT 100.340 136.570 261.550 136.620 ;
        RECT 98.750 136.100 261.550 136.570 ;
        RECT 98.750 136.050 100.670 136.100 ;
        RECT 98.750 121.475 99.270 136.050 ;
        RECT 98.745 120.945 99.275 121.475 ;
        RECT 101.335 119.960 130.945 134.505 ;
        RECT 132.935 119.960 162.545 134.505 ;
        RECT 164.535 119.960 194.145 134.505 ;
        RECT 196.135 119.960 225.745 134.505 ;
        RECT 227.735 119.960 257.345 134.505 ;
        RECT 258.150 119.960 260.190 120.020 ;
        RECT 96.610 119.500 260.190 119.960 ;
        RECT 96.610 119.440 258.340 119.500 ;
        RECT -323.040 118.380 59.490 118.450 ;
        RECT -323.040 117.930 63.040 118.380 ;
        RECT -321.130 102.050 -320.610 117.160 ;
        RECT -318.715 103.385 -289.105 117.930 ;
        RECT -287.115 103.385 -257.505 117.930 ;
        RECT -255.515 103.385 -225.905 117.930 ;
        RECT -223.915 103.385 -194.305 117.930 ;
        RECT -192.315 103.385 -162.705 117.930 ;
        RECT -160.715 103.385 -131.105 117.930 ;
        RECT -129.115 103.385 -99.505 117.930 ;
        RECT -97.515 103.385 -67.905 117.930 ;
        RECT -65.915 103.385 -36.305 117.930 ;
        RECT -34.315 103.385 -4.705 117.930 ;
        RECT -2.715 103.385 26.895 117.930 ;
        RECT 28.885 103.385 58.495 117.930 ;
        RECT 59.140 117.860 63.040 117.930 ;
        RECT 59.040 102.050 60.750 102.140 ;
        RECT -321.130 101.620 60.750 102.050 ;
        RECT -321.130 101.530 59.490 101.620 ;
        RECT -318.715 85.390 -289.105 99.935 ;
        RECT -287.115 85.390 -257.505 99.935 ;
        RECT -255.515 85.390 -225.905 99.935 ;
        RECT -223.915 85.390 -194.305 99.935 ;
        RECT -192.315 85.390 -162.705 99.935 ;
        RECT -160.715 85.390 -131.105 99.935 ;
        RECT -129.115 85.390 -99.505 99.935 ;
        RECT -97.515 85.390 -67.905 99.935 ;
        RECT -65.915 85.390 -36.305 99.935 ;
        RECT -34.315 85.390 -4.705 99.935 ;
        RECT -2.715 85.390 26.895 99.935 ;
        RECT 28.885 85.390 58.495 99.935 ;
        RECT 60.230 86.445 60.750 101.620 ;
        RECT 60.225 85.915 60.755 86.445 ;
        RECT 62.520 85.390 63.040 117.860 ;
        RECT 98.750 103.560 99.270 118.400 ;
        RECT 101.335 104.895 130.945 119.440 ;
        RECT 132.935 104.895 162.545 119.440 ;
        RECT 164.535 104.895 194.145 119.440 ;
        RECT 196.135 104.895 225.745 119.440 ;
        RECT 227.735 104.895 257.345 119.440 ;
        RECT 258.735 103.580 259.265 103.585 ;
        RECT 257.790 103.560 259.265 103.580 ;
        RECT 98.750 103.060 259.265 103.560 ;
        RECT 98.750 103.040 258.340 103.060 ;
        RECT 258.735 103.055 259.265 103.060 ;
        RECT 101.335 86.900 130.945 101.445 ;
        RECT 132.935 86.900 162.545 101.445 ;
        RECT 164.535 86.900 194.145 101.445 ;
        RECT 196.135 86.900 225.745 101.445 ;
        RECT 227.735 86.900 257.345 101.445 ;
        RECT 259.670 86.900 260.190 119.500 ;
        RECT 91.525 86.880 91.975 86.885 ;
        RECT 100.340 86.880 260.190 86.900 ;
        RECT 91.525 86.440 260.190 86.880 ;
        RECT 91.525 86.435 91.975 86.440 ;
        RECT 100.340 86.380 260.190 86.440 ;
        RECT -319.710 85.240 63.040 85.390 ;
        RECT -323.830 84.870 63.040 85.240 ;
        RECT -323.830 84.720 -319.240 84.870 ;
        RECT -323.830 52.330 -323.310 84.720 ;
        RECT -318.715 70.325 -289.105 84.870 ;
        RECT -287.115 70.325 -257.505 84.870 ;
        RECT -255.515 70.325 -225.905 84.870 ;
        RECT -223.915 70.325 -194.305 84.870 ;
        RECT -192.315 70.325 -162.705 84.870 ;
        RECT -160.715 70.325 -131.105 84.870 ;
        RECT -129.115 70.325 -99.505 84.870 ;
        RECT -97.515 70.325 -67.905 84.870 ;
        RECT -65.915 70.325 -36.305 84.870 ;
        RECT -34.315 70.325 -4.705 84.870 ;
        RECT -2.715 70.325 26.895 84.870 ;
        RECT 28.885 70.325 58.495 84.870 ;
        RECT -322.000 68.990 -319.080 69.040 ;
        RECT 60.230 68.990 60.750 84.120 ;
        RECT 86.025 76.120 86.555 76.125 ;
        RECT 86.025 75.600 99.240 76.120 ;
        RECT 86.025 75.595 86.555 75.600 ;
        RECT 98.720 70.480 99.240 75.600 ;
        RECT 101.335 71.835 130.945 86.380 ;
        RECT 132.935 71.835 162.545 86.380 ;
        RECT 164.535 71.835 194.145 86.380 ;
        RECT 196.135 71.835 225.745 86.380 ;
        RECT 227.735 71.835 257.345 86.380 ;
        RECT 261.400 70.500 261.920 103.580 ;
        RECT 100.340 70.480 261.920 70.500 ;
        RECT 98.720 69.980 261.920 70.480 ;
        RECT 98.720 69.960 100.790 69.980 ;
        RECT -322.000 68.520 60.750 68.990 ;
        RECT -322.000 54.395 -321.480 68.520 ;
        RECT -319.710 68.470 60.750 68.520 ;
        RECT -322.005 53.865 -321.475 54.395 ;
        RECT -318.715 52.330 -289.105 66.875 ;
        RECT -287.115 52.330 -257.505 66.875 ;
        RECT -255.515 52.330 -225.905 66.875 ;
        RECT -223.915 52.330 -194.305 66.875 ;
        RECT -192.315 52.330 -162.705 66.875 ;
        RECT -160.715 52.330 -131.105 66.875 ;
        RECT -129.115 52.330 -99.505 66.875 ;
        RECT -97.515 52.330 -67.905 66.875 ;
        RECT -65.915 52.330 -36.305 66.875 ;
        RECT -34.315 52.330 -4.705 66.875 ;
        RECT -2.715 52.330 26.895 66.875 ;
        RECT 28.885 52.330 58.495 66.875 ;
        RECT -323.830 51.810 60.770 52.330 ;
        RECT -322.000 35.930 -321.480 50.820 ;
        RECT -318.715 37.265 -289.105 51.810 ;
        RECT -287.115 37.265 -257.505 51.810 ;
        RECT -255.515 37.265 -225.905 51.810 ;
        RECT -223.915 37.265 -194.305 51.810 ;
        RECT -192.315 37.265 -162.705 51.810 ;
        RECT -160.715 37.265 -131.105 51.810 ;
        RECT -129.115 37.265 -99.505 51.810 ;
        RECT -97.515 37.265 -67.905 51.810 ;
        RECT -65.915 37.265 -36.305 51.810 ;
        RECT -34.315 37.265 -4.705 51.810 ;
        RECT -2.715 37.265 26.895 51.810 ;
        RECT 28.885 37.265 58.495 51.810 ;
        RECT -322.000 35.900 60.510 35.930 ;
        RECT 63.025 35.900 63.555 35.905 ;
        RECT -322.000 35.410 63.555 35.900 ;
        RECT 59.940 35.380 63.555 35.410 ;
        RECT 63.025 35.375 63.555 35.380 ;
  END
END pll
END LIBRARY

