# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nor4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 2.275000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.995000 1.785000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.995000 1.285000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.795000 1.615000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.871000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.655000 1.925000 0.825000 ;
        RECT 0.085000 0.825000 0.345000 2.450000 ;
        RECT 0.855000 0.300000 1.055000 0.655000 ;
        RECT 1.725000 0.310000 1.925000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.355000  0.085000 0.685000 0.480000 ;
        RECT 1.225000  0.085000 1.555000 0.485000 ;
        RECT 2.095000  0.085000 2.425000 0.825000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 2.095000 2.185000 2.425000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525000 0.995000 0.745000 1.795000 ;
      RECT 0.525000 1.795000 3.135000 2.005000 ;
      RECT 2.660000 0.405000 2.830000 0.655000 ;
      RECT 2.660000 0.655000 3.135000 0.825000 ;
      RECT 2.965000 0.825000 3.135000 1.795000 ;
  END
END sky130_fd_sc_hd__nor4b_1
END LIBRARY
