# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__or3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 1.075000 2.230000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 2.125000 3.135000 2.365000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.265000 1.285000 0.595000 ;
        RECT 0.935000 0.595000 1.105000 1.495000 ;
        RECT 0.935000 1.495000 1.330000 1.700000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.595000  0.085000 0.765000 0.565000 ;
        RECT 1.520000  0.085000 1.690000 0.565000 ;
        RECT 2.330000  0.085000 2.660000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.550000 2.210000 0.910000 2.635000 ;
        RECT 1.425000 2.210000 1.755000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.290000 0.345000 0.735000 ;
      RECT 0.085000 0.735000 0.765000 0.905000 ;
      RECT 0.085000 1.810000 0.765000 1.870000 ;
      RECT 0.085000 1.870000 2.660000 1.955000 ;
      RECT 0.085000 1.955000 1.720000 2.040000 ;
      RECT 0.085000 2.040000 0.345000 2.220000 ;
      RECT 0.595000 0.905000 0.765000 1.810000 ;
      RECT 1.275000 0.765000 3.135000 0.825000 ;
      RECT 1.275000 0.825000 2.160000 0.905000 ;
      RECT 1.275000 0.905000 1.595000 0.935000 ;
      RECT 1.275000 0.935000 1.445000 1.325000 ;
      RECT 1.425000 0.735000 3.135000 0.765000 ;
      RECT 1.550000 1.785000 2.660000 1.870000 ;
      RECT 1.990000 0.305000 2.160000 0.655000 ;
      RECT 1.990000 0.655000 3.135000 0.735000 ;
      RECT 2.490000 0.995000 2.790000 1.325000 ;
      RECT 2.490000 1.325000 2.660000 1.785000 ;
      RECT 2.830000 0.305000 3.085000 0.605000 ;
      RECT 2.830000 0.605000 3.135000 0.655000 ;
      RECT 2.830000 1.495000 3.135000 1.925000 ;
      RECT 2.965000 0.825000 3.135000 1.495000 ;
  END
END sky130_fd_sc_hd__or3b_2
END LIBRARY
