# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a21boi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 1.065000 4.970000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.030000 1.065000 3.375000 1.480000 ;
        RECT 3.030000 1.480000 6.450000 1.705000 ;
        RECT 5.205000 1.075000 6.450000 1.480000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.650000 1.615000 ;
        RECT 0.480000 0.995000 0.650000 1.075000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 0.370000 1.465000 0.615000 ;
        RECT 1.275000 0.615000 2.325000 0.695000 ;
        RECT 1.275000 0.695000 4.885000 0.865000 ;
        RECT 1.560000 1.585000 2.860000 1.705000 ;
        RECT 1.560000 1.705000 2.725000 2.035000 ;
        RECT 2.135000 0.255000 2.325000 0.615000 ;
        RECT 2.570000 0.865000 4.885000 0.895000 ;
        RECT 2.570000 0.895000 2.860000 1.585000 ;
        RECT 3.255000 0.675000 4.885000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.720000  0.085000 1.105000 0.445000 ;
        RECT 1.635000  0.085000 1.965000 0.445000 ;
        RECT 2.495000  0.085000 3.085000 0.525000 ;
        RECT 5.485000  0.085000 5.675000 0.565000 ;
        RECT 6.345000  0.085000 6.605000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.625000 2.175000 0.885000 2.635000 ;
        RECT 3.265000 2.275000 3.595000 2.635000 ;
        RECT 4.125000 2.275000 4.455000 2.635000 ;
        RECT 4.985000 2.275000 5.315000 2.635000 ;
        RECT 5.845000 2.275000 6.175000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.445000 0.615000 ;
      RECT 0.090000 0.615000 1.105000 0.795000 ;
      RECT 0.125000 1.785000 0.990000 2.005000 ;
      RECT 0.125000 2.005000 0.455000 2.465000 ;
      RECT 0.820000 0.795000 1.105000 1.035000 ;
      RECT 0.820000 1.035000 2.400000 1.345000 ;
      RECT 0.820000 1.345000 0.990000 1.785000 ;
      RECT 1.160000 1.795000 1.355000 2.215000 ;
      RECT 1.160000 2.215000 3.095000 2.465000 ;
      RECT 1.935000 2.205000 3.095000 2.215000 ;
      RECT 2.895000 1.875000 6.605000 2.105000 ;
      RECT 2.895000 2.105000 3.095000 2.205000 ;
      RECT 3.265000 0.255000 5.315000 0.505000 ;
      RECT 4.625000 2.105000 4.815000 2.465000 ;
      RECT 5.055000 0.505000 5.315000 0.735000 ;
      RECT 5.055000 0.735000 6.175000 0.905000 ;
      RECT 5.485000 2.105000 5.665000 2.465000 ;
      RECT 5.845000 0.255000 6.175000 0.735000 ;
      RECT 6.345000 2.105000 6.605000 2.465000 ;
  END
END sky130_fd_sc_hd__a21boi_4
END LIBRARY
