# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.110000 0.795000 ;
        RECT 8.855000 1.445000 9.110000 2.325000 ;
        RECT 8.900000 0.795000 9.110000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.200000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.465000 ;
        RECT 1.545000  0.085000 1.875000 0.445000 ;
        RECT 4.475000  0.085000 4.805000 0.545000 ;
        RECT 6.705000  0.085000 6.895000 0.525000 ;
        RECT 8.380000  0.085000 8.685000 0.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.200000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.850000 2.175000 2.100000 2.635000 ;
        RECT 3.990000 2.205000 4.320000 2.635000 ;
        RECT 4.955000 2.175000 5.325000 2.635000 ;
        RECT 6.940000 2.175000 7.190000 2.635000 ;
        RECT 7.710000 2.255000 8.040000 2.635000 ;
        RECT 8.380000 1.495000 8.685000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.345000 0.345000 0.635000 ;
      RECT 0.090000 0.635000 0.840000 0.805000 ;
      RECT 0.090000 1.795000 0.840000 1.965000 ;
      RECT 0.090000 1.965000 0.345000 2.465000 ;
      RECT 0.610000 0.805000 0.840000 1.795000 ;
      RECT 1.015000 0.345000 1.185000 2.465000 ;
      RECT 2.045000 0.305000 2.540000 0.475000 ;
      RECT 2.045000 0.475000 2.215000 1.835000 ;
      RECT 2.045000 1.835000 2.440000 2.005000 ;
      RECT 2.270000 2.005000 2.440000 2.135000 ;
      RECT 2.270000 2.135000 2.520000 2.465000 ;
      RECT 2.385000 0.765000 2.735000 1.385000 ;
      RECT 2.610000 1.575000 3.075000 1.965000 ;
      RECT 2.735000 2.135000 3.415000 2.465000 ;
      RECT 2.745000 0.305000 3.600000 0.475000 ;
      RECT 2.905000 0.765000 3.260000 0.985000 ;
      RECT 2.905000 0.985000 3.075000 1.575000 ;
      RECT 3.245000 1.185000 4.935000 1.355000 ;
      RECT 3.245000 1.355000 3.415000 2.135000 ;
      RECT 3.430000 0.475000 3.600000 1.185000 ;
      RECT 3.585000 1.865000 4.660000 2.035000 ;
      RECT 3.585000 2.035000 3.755000 2.375000 ;
      RECT 3.775000 1.525000 5.275000 1.695000 ;
      RECT 4.490000 2.035000 4.660000 2.375000 ;
      RECT 4.765000 1.005000 4.935000 1.185000 ;
      RECT 5.015000 0.275000 5.365000 0.445000 ;
      RECT 5.015000 0.445000 5.275000 0.835000 ;
      RECT 5.105000 0.835000 5.275000 1.525000 ;
      RECT 5.105000 1.695000 5.275000 1.835000 ;
      RECT 5.105000 1.835000 5.665000 2.005000 ;
      RECT 5.465000 0.705000 5.675000 1.495000 ;
      RECT 5.465000 1.495000 6.140000 1.655000 ;
      RECT 5.465000 1.655000 6.430000 1.665000 ;
      RECT 5.495000 2.005000 5.665000 2.465000 ;
      RECT 5.585000 0.255000 6.535000 0.535000 ;
      RECT 5.845000 0.705000 6.195000 1.325000 ;
      RECT 5.900000 2.125000 6.770000 2.465000 ;
      RECT 5.970000 1.665000 6.430000 1.955000 ;
      RECT 6.365000 0.535000 6.535000 1.315000 ;
      RECT 6.365000 1.315000 6.770000 1.485000 ;
      RECT 6.600000 1.485000 6.770000 1.575000 ;
      RECT 6.600000 1.575000 7.820000 1.745000 ;
      RECT 6.600000 1.745000 6.770000 2.125000 ;
      RECT 6.705000 0.695000 7.235000 0.865000 ;
      RECT 6.705000 0.865000 6.925000 1.145000 ;
      RECT 7.065000 0.295000 8.135000 0.465000 ;
      RECT 7.065000 0.465000 7.235000 0.695000 ;
      RECT 7.360000 1.915000 8.160000 2.085000 ;
      RECT 7.360000 2.085000 7.530000 2.375000 ;
      RECT 7.815000 0.465000 8.135000 0.820000 ;
      RECT 7.815000 0.820000 8.140000 0.995000 ;
      RECT 7.815000 0.995000 8.730000 1.295000 ;
      RECT 7.990000 1.295000 8.730000 1.325000 ;
      RECT 7.990000 1.325000 8.160000 1.915000 ;
    LAYER mcon ;
      RECT 0.610000 1.105000 0.780000 1.275000 ;
      RECT 1.015000 1.785000 1.185000 1.955000 ;
      RECT 2.445000 1.105000 2.615000 1.275000 ;
      RECT 2.905000 1.785000 3.075000 1.955000 ;
      RECT 6.025000 1.105000 6.195000 1.275000 ;
      RECT 6.025000 1.785000 6.195000 1.955000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_1
END LIBRARY
