# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o311a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.950000 1.055000 7.735000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.020000 1.055000 6.770000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 1.055000 5.850000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.055000 4.475000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.115000 1.055000 3.080000 1.315000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.765000 1.315000 ;
        RECT 0.595000 0.255000 0.765000 0.715000 ;
        RECT 0.595000 0.715000 1.605000 0.885000 ;
        RECT 0.595000 0.885000 0.765000 1.055000 ;
        RECT 0.595000 1.315000 0.765000 1.485000 ;
        RECT 0.595000 1.485000 1.605000 1.725000 ;
        RECT 0.595000 1.725000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.715000 ;
        RECT 1.435000 1.725000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.085000  0.085000 0.425000 0.885000 ;
        RECT 0.935000  0.085000 1.265000 0.545000 ;
        RECT 1.775000  0.085000 2.025000 0.545000 ;
        RECT 4.925000  0.085000 5.605000 0.505000 ;
        RECT 6.115000  0.085000 6.445000 0.505000 ;
        RECT 6.955000  0.085000 7.285000 0.505000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.085000 1.485000 0.425000 2.635000 ;
        RECT 0.935000 1.895000 1.265000 2.635000 ;
        RECT 1.775000 1.895000 2.445000 2.635000 ;
        RECT 2.955000 1.895000 3.285000 2.635000 ;
        RECT 3.855000 1.895000 4.045000 2.635000 ;
        RECT 6.955000 1.895000 7.285000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.935000 1.055000 1.945000 1.315000 ;
      RECT 1.775000 0.715000 3.045000 0.885000 ;
      RECT 1.775000 0.885000 1.945000 1.055000 ;
      RECT 1.775000 1.315000 1.945000 1.485000 ;
      RECT 1.775000 1.485000 5.005000 1.725000 ;
      RECT 2.195000 0.255000 4.305000 0.505000 ;
      RECT 2.195000 0.675000 3.045000 0.715000 ;
      RECT 2.615000 1.725000 2.785000 2.465000 ;
      RECT 3.215000 0.505000 3.385000 0.885000 ;
      RECT 3.455000 1.725000 3.625000 2.465000 ;
      RECT 3.555000 0.675000 7.735000 0.885000 ;
      RECT 4.335000 1.895000 4.665000 2.295000 ;
      RECT 4.335000 2.295000 6.445000 2.465000 ;
      RECT 4.485000 0.255000 4.755000 0.675000 ;
      RECT 4.835000 1.725000 5.005000 2.125000 ;
      RECT 5.255000 1.485000 5.525000 2.295000 ;
      RECT 5.695000 1.485000 7.735000 1.725000 ;
      RECT 5.695000 1.725000 5.945000 2.125000 ;
      RECT 5.775000 0.255000 5.945000 0.675000 ;
      RECT 6.115000 1.895000 6.445000 2.295000 ;
      RECT 6.615000 0.255000 6.785000 0.675000 ;
      RECT 6.615000 1.725000 6.785000 2.125000 ;
      RECT 7.455000 0.255000 7.735000 0.675000 ;
      RECT 7.455000 1.725000 7.735000 2.465000 ;
  END
END sky130_fd_sc_hd__o311a_4
END LIBRARY
