# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__fahcin_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.665000 1.740000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.240000 0.645000 4.490000 1.325000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 0.735000 1.755000 0.780000 ;
        RECT 1.465000 0.780000 4.515000 0.920000 ;
        RECT 1.465000 0.920000 1.755000 0.965000 ;
        RECT 4.225000 0.735000 4.515000 0.780000 ;
        RECT 4.225000 0.920000 4.515000 0.965000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.520000 1.075000 10.965000 1.275000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.600000 0.755000 6.925000 0.925000 ;
        RECT 6.600000 0.925000 6.870000 1.675000 ;
        RECT 6.700000 1.675000 6.870000 1.785000 ;
        RECT 6.755000 0.595000 6.925000 0.755000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.255000 12.335000 0.825000 ;
        RECT 12.000000 1.785000 12.335000 2.465000 ;
        RECT 12.125000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.420000 0.085000 ;
        RECT  0.630000  0.085000  0.800000 0.545000 ;
        RECT  5.180000  0.085000  5.510000 0.805000 ;
        RECT 10.180000  0.085000 10.350000 0.565000 ;
        RECT 11.495000  0.085000 11.825000 0.510000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 12.420000 2.805000 ;
        RECT  0.600000 2.180000  0.770000 2.635000 ;
        RECT  5.260000 2.235000  5.590000 2.635000 ;
        RECT 10.190000 2.195000 10.360000 2.635000 ;
        RECT 11.575000 1.785000 11.830000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.735000  0.430000 0.805000 ;
      RECT  0.085000 0.805000  0.255000 1.500000 ;
      RECT  0.085000 1.500000  0.440000 1.840000 ;
      RECT  0.085000 1.840000  1.110000 2.010000 ;
      RECT  0.085000 2.010000  0.430000 2.465000 ;
      RECT  0.100000 0.255000  0.430000 0.735000 ;
      RECT  0.425000 0.995000  0.780000 1.325000 ;
      RECT  0.610000 0.735000  1.325000 0.905000 ;
      RECT  0.610000 0.905000  0.780000 0.995000 ;
      RECT  0.610000 1.325000  0.780000 1.500000 ;
      RECT  0.610000 1.500000  1.450000 1.670000 ;
      RECT  0.940000 2.010000  1.110000 2.215000 ;
      RECT  0.940000 2.215000  1.970000 2.295000 ;
      RECT  0.940000 2.295000  3.515000 2.385000 ;
      RECT  0.995000 0.255000  3.390000 0.425000 ;
      RECT  0.995000 0.425000  2.100000 0.465000 ;
      RECT  0.995000 0.465000  1.325000 0.735000 ;
      RECT  1.280000 1.670000  1.450000 1.785000 ;
      RECT  1.280000 1.785000  2.050000 1.955000 ;
      RECT  1.280000 1.955000  1.450000 2.045000 ;
      RECT  1.715000 2.385000  3.515000 2.465000 ;
      RECT  1.985000 0.675000  2.390000 1.350000 ;
      RECT  2.220000 0.595000  2.390000 0.675000 ;
      RECT  2.220000 1.350000  2.390000 1.785000 ;
      RECT  2.515000 0.425000  3.390000 0.465000 ;
      RECT  2.565000 1.785000  2.895000 2.045000 ;
      RECT  2.620000 0.655000  3.025000 0.735000 ;
      RECT  2.620000 0.735000  3.135000 0.755000 ;
      RECT  2.620000 0.755000  3.730000 0.905000 ;
      RECT  2.640000 1.075000  2.970000 1.095000 ;
      RECT  2.640000 1.095000  3.120000 1.245000 ;
      RECT  2.800000 1.245000  3.120000 1.265000 ;
      RECT  2.950000 1.265000  3.120000 1.615000 ;
      RECT  3.055000 0.905000  3.730000 0.925000 ;
      RECT  3.215000 0.465000  3.390000 0.585000 ;
      RECT  3.245000 2.110000  3.460000 2.295000 ;
      RECT  3.290000 0.925000  3.460000 2.110000 ;
      RECT  3.560000 0.255000  4.570000 0.425000 ;
      RECT  3.560000 0.425000  3.730000 0.755000 ;
      RECT  3.710000 1.150000  4.070000 1.320000 ;
      RECT  3.710000 1.320000  3.880000 2.290000 ;
      RECT  3.710000 2.290000  5.065000 2.460000 ;
      RECT  3.900000 0.595000  4.070000 1.150000 ;
      RECT  4.080000 1.695000  4.445000 2.120000 ;
      RECT  4.240000 0.425000  4.570000 0.475000 ;
      RECT  4.690000 1.385000  5.170000 1.725000 ;
      RECT  4.815000 1.895000  5.995000 2.065000 ;
      RECT  4.815000 2.065000  5.065000 2.290000 ;
      RECT  4.830000 0.510000  5.000000 0.995000 ;
      RECT  4.830000 0.995000  5.630000 1.325000 ;
      RECT  4.830000 1.325000  5.170000 1.385000 ;
      RECT  5.635000 1.555000  6.370000 1.725000 ;
      RECT  5.680000 0.380000  5.970000 0.815000 ;
      RECT  5.800000 0.815000  5.970000 1.555000 ;
      RECT  5.825000 2.065000  5.995000 2.295000 ;
      RECT  5.825000 2.295000  7.950000 2.465000 ;
      RECT  6.140000 0.740000  6.425000 1.325000 ;
      RECT  6.200000 1.725000  6.370000 1.895000 ;
      RECT  6.200000 1.895000  6.530000 1.955000 ;
      RECT  6.200000 1.955000  7.210000 2.125000 ;
      RECT  6.255000 0.255000  7.695000 0.425000 ;
      RECT  6.255000 0.425000  6.585000 0.570000 ;
      RECT  7.040000 1.060000  7.270000 1.230000 ;
      RECT  7.040000 1.230000  7.210000 1.955000 ;
      RECT  7.100000 0.595000  7.350000 0.925000 ;
      RECT  7.100000 0.925000  7.270000 1.060000 ;
      RECT  7.380000 1.360000  7.610000 1.530000 ;
      RECT  7.380000 1.530000  7.550000 2.125000 ;
      RECT  7.440000 1.105000  7.695000 1.290000 ;
      RECT  7.440000 1.290000  7.610000 1.360000 ;
      RECT  7.520000 0.425000  7.695000 1.105000 ;
      RECT  7.780000 1.550000  8.035000 1.720000 ;
      RECT  7.780000 1.720000  7.950000 2.295000 ;
      RECT  7.865000 0.255000  9.980000 0.425000 ;
      RECT  7.865000 0.425000  8.035000 0.740000 ;
      RECT  7.865000 0.995000  8.035000 1.550000 ;
      RECT  8.220000 1.955000  8.390000 2.295000 ;
      RECT  8.220000 2.295000  9.410000 2.465000 ;
      RECT  8.305000 0.595000  8.555000 0.925000 ;
      RECT  8.375000 0.925000  8.555000 1.445000 ;
      RECT  8.375000 1.445000  8.670000 1.530000 ;
      RECT  8.375000 1.530000  8.890000 1.785000 ;
      RECT  8.560000 1.785000  8.890000 2.125000 ;
      RECT  8.725000 0.595000  9.410000 0.765000 ;
      RECT  8.835000 0.995000  9.070000 1.325000 ;
      RECT  9.240000 0.765000  9.410000 1.875000 ;
      RECT  9.240000 1.875000 10.885000 2.025000 ;
      RECT  9.240000 2.025000 10.145000 2.030000 ;
      RECT  9.240000 2.030000 10.130000 2.035000 ;
      RECT  9.240000 2.035000 10.120000 2.040000 ;
      RECT  9.240000 2.040000 10.105000 2.045000 ;
      RECT  9.240000 2.045000  9.410000 2.295000 ;
      RECT  9.640000 0.425000  9.980000 0.825000 ;
      RECT  9.640000 0.825000  9.810000 1.535000 ;
      RECT  9.640000 1.535000 10.010000 1.705000 ;
      RECT  9.980000 0.995000 10.350000 1.325000 ;
      RECT 10.055000 1.870000 10.885000 1.875000 ;
      RECT 10.070000 1.865000 10.885000 1.870000 ;
      RECT 10.085000 1.860000 10.885000 1.865000 ;
      RECT 10.100000 1.855000 10.885000 1.860000 ;
      RECT 10.180000 0.735000 10.910000 0.905000 ;
      RECT 10.180000 0.905000 10.350000 0.995000 ;
      RECT 10.180000 1.325000 10.350000 1.445000 ;
      RECT 10.180000 1.445000 10.885000 1.855000 ;
      RECT 10.530000 0.285000 10.910000 0.735000 ;
      RECT 10.535000 2.025000 10.885000 2.465000 ;
      RECT 11.075000 1.455000 11.405000 2.465000 ;
      RECT 11.155000 0.270000 11.325000 0.680000 ;
      RECT 11.155000 0.680000 11.405000 1.455000 ;
      RECT 11.645000 0.995000 11.955000 1.615000 ;
    LAYER mcon ;
      RECT  1.880000 1.785000  2.050000 1.955000 ;
      RECT  1.985000 1.105000  2.155000 1.275000 ;
      RECT  2.570000 1.785000  2.740000 1.955000 ;
      RECT  2.950000 1.445000  3.120000 1.615000 ;
      RECT  4.140000 1.785000  4.310000 1.955000 ;
      RECT  4.760000 1.445000  4.930000 1.615000 ;
      RECT  6.140000 1.105000  6.310000 1.275000 ;
      RECT  7.520000 0.765000  7.690000 0.935000 ;
      RECT  8.440000 1.445000  8.610000 1.615000 ;
      RECT  8.900000 1.105000  9.070000 1.275000 ;
      RECT 11.220000 0.765000 11.390000 0.935000 ;
      RECT 11.680000 1.445000 11.850000 1.615000 ;
    LAYER met1 ;
      RECT  1.820000 1.755000  2.110000 1.800000 ;
      RECT  1.820000 1.800000  4.370000 1.940000 ;
      RECT  1.820000 1.940000  2.110000 1.985000 ;
      RECT  1.925000 1.075000  2.215000 1.120000 ;
      RECT  1.925000 1.120000  9.130000 1.260000 ;
      RECT  1.925000 1.260000  2.215000 1.305000 ;
      RECT  2.510000 1.755000  2.800000 1.800000 ;
      RECT  2.510000 1.940000  2.800000 1.985000 ;
      RECT  2.890000 1.415000  3.180000 1.460000 ;
      RECT  2.890000 1.460000  4.990000 1.600000 ;
      RECT  2.890000 1.600000  3.180000 1.645000 ;
      RECT  4.080000 1.755000  4.370000 1.800000 ;
      RECT  4.080000 1.940000  4.370000 1.985000 ;
      RECT  4.700000 1.415000  4.990000 1.460000 ;
      RECT  4.700000 1.600000  4.990000 1.645000 ;
      RECT  6.080000 1.075000  6.370000 1.120000 ;
      RECT  6.080000 1.260000  6.370000 1.305000 ;
      RECT  7.460000 0.735000  7.750000 0.780000 ;
      RECT  7.460000 0.780000 11.450000 0.920000 ;
      RECT  7.460000 0.920000  7.750000 0.965000 ;
      RECT  8.380000 1.415000  8.670000 1.460000 ;
      RECT  8.380000 1.460000 11.910000 1.600000 ;
      RECT  8.380000 1.600000  8.670000 1.645000 ;
      RECT  8.840000 1.075000  9.130000 1.120000 ;
      RECT  8.840000 1.260000  9.130000 1.305000 ;
      RECT 11.160000 0.735000 11.450000 0.780000 ;
      RECT 11.160000 0.920000 11.450000 0.965000 ;
      RECT 11.620000 1.415000 11.910000 1.460000 ;
      RECT 11.620000 1.600000 11.910000 1.645000 ;
  END
END sky130_fd_sc_hd__fahcin_1
END LIBRARY
