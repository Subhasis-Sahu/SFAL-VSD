# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__fa_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 0.995000 1.755000 1.275000 ;
        RECT 1.245000 1.275000 1.505000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685000 1.030000 3.075000 1.360000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.720000 0.955000 5.080000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.105000 0.995000 6.960000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000 1.755000 1.120000 ;
        RECT 1.465000 1.120000 6.375000 1.260000 ;
        RECT 1.465000 1.260000 1.755000 1.305000 ;
        RECT 2.845000 1.075000 3.135000 1.120000 ;
        RECT 2.845000 1.260000 3.135000 1.305000 ;
        RECT 4.705000 1.075000 4.995000 1.120000 ;
        RECT 4.705000 1.260000 4.995000 1.305000 ;
        RECT 6.085000 1.075000 6.375000 1.120000 ;
        RECT 6.085000 1.260000 6.375000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645000 1.445000 2.155000 1.690000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.655000 1.435000 4.070000 1.745000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.150000 1.445000 6.835000 1.735000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.925000 1.415000 2.215000 1.460000 ;
        RECT 1.925000 1.460000 6.835000 1.600000 ;
        RECT 1.925000 1.600000 2.215000 1.645000 ;
        RECT 3.785000 1.415000 4.075000 1.460000 ;
        RECT 3.785000 1.600000 4.075000 1.645000 ;
        RECT 6.545000 1.415000 6.835000 1.460000 ;
        RECT 6.545000 1.600000 6.835000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.475500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 1.105000 2.495000 1.275000 ;
        RECT 2.325000 1.275000 2.495000 1.570000 ;
        RECT 2.325000 1.570000 3.415000 1.740000 ;
        RECT 3.245000 0.965000 4.465000 1.250000 ;
        RECT 3.245000 1.250000 3.415000 1.570000 ;
        RECT 4.295000 1.250000 4.465000 1.435000 ;
        RECT 4.295000 1.435000 4.655000 1.515000 ;
        RECT 4.295000 1.515000 5.920000 1.685000 ;
        RECT 5.670000 1.355000 5.920000 1.515000 ;
        RECT 5.670000 1.685000 5.920000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.735000 0.690000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.415000 ;
        RECT 0.085000 1.415000 0.735000 1.585000 ;
        RECT 0.520000 0.315000 0.850000 0.485000 ;
        RECT 0.520000 0.485000 0.690000 0.735000 ;
        RECT 0.565000 1.585000 0.735000 1.780000 ;
        RECT 0.565000 1.780000 0.810000 1.950000 ;
        RECT 0.600000 1.950000 0.810000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.523500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.395000 0.255000 7.725000 0.485000 ;
        RECT 7.395000 1.795000 7.645000 1.965000 ;
        RECT 7.395000 1.965000 7.565000 2.465000 ;
        RECT 7.475000 0.485000 7.725000 0.735000 ;
        RECT 7.475000 0.735000 8.195000 0.905000 ;
        RECT 7.475000 1.415000 8.195000 1.585000 ;
        RECT 7.475000 1.585000 7.645000 1.795000 ;
        RECT 7.970000 0.905000 8.195000 1.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 0.180000  0.085000 0.350000 0.565000 ;
        RECT 1.020000  0.085000 1.350000 0.465000 ;
        RECT 2.755000  0.085000 3.085000 0.445000 ;
        RECT 3.695000  0.085000 4.025000 0.490000 ;
        RECT 4.535000  0.085000 4.865000 0.445000 ;
        RECT 6.780000  0.085000 7.110000 0.445000 ;
        RECT 7.895000  0.085000 8.065000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 0.180000 1.795000 0.350000 2.635000 ;
        RECT 0.980000 2.275000 1.310000 2.635000 ;
        RECT 2.755000 2.275000 3.085000 2.635000 ;
        RECT 3.695000 1.915000 4.025000 2.635000 ;
        RECT 4.535000 2.275000 4.865000 2.635000 ;
        RECT 6.890000 2.275000 7.220000 2.635000 ;
        RECT 7.815000 1.795000 7.985000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.540000 1.075000 1.075000 1.245000 ;
      RECT 0.905000 0.655000 2.165000 0.825000 ;
      RECT 0.905000 0.825000 1.075000 1.075000 ;
      RECT 0.905000 1.245000 1.075000 1.430000 ;
      RECT 0.905000 1.430000 1.110000 1.495000 ;
      RECT 0.905000 1.495000 1.475000 1.600000 ;
      RECT 0.940000 1.600000 1.475000 1.665000 ;
      RECT 1.305000 1.665000 1.475000 1.910000 ;
      RECT 1.305000 1.910000 2.245000 2.080000 ;
      RECT 1.535000 0.255000 2.165000 0.655000 ;
      RECT 1.900000 2.080000 2.245000 2.465000 ;
      RECT 1.925000 0.825000 2.165000 0.935000 ;
      RECT 2.415000 0.255000 2.585000 0.615000 ;
      RECT 2.415000 0.615000 3.425000 0.785000 ;
      RECT 2.415000 1.935000 3.490000 2.105000 ;
      RECT 2.415000 2.105000 2.585000 2.465000 ;
      RECT 3.255000 0.255000 3.425000 0.615000 ;
      RECT 3.255000 2.105000 3.490000 2.465000 ;
      RECT 4.195000 0.255000 4.365000 0.615000 ;
      RECT 4.195000 0.615000 5.205000 0.785000 ;
      RECT 4.195000 1.935000 5.205000 2.105000 ;
      RECT 4.195000 2.105000 4.365000 2.465000 ;
      RECT 5.035000 0.255000 5.205000 0.615000 ;
      RECT 5.035000 2.105000 5.205000 2.465000 ;
      RECT 5.250000 0.955000 5.935000 1.125000 ;
      RECT 5.420000 0.765000 5.935000 0.955000 ;
      RECT 5.485000 2.125000 6.685000 2.465000 ;
      RECT 5.540000 0.255000 6.550000 0.505000 ;
      RECT 5.540000 0.505000 5.710000 0.595000 ;
      RECT 6.380000 0.505000 6.550000 0.655000 ;
      RECT 6.380000 0.655000 7.300000 0.825000 ;
      RECT 6.515000 1.935000 7.180000 2.105000 ;
      RECT 6.515000 2.105000 6.685000 2.125000 ;
      RECT 7.010000 1.470000 7.300000 1.640000 ;
      RECT 7.010000 1.640000 7.180000 1.935000 ;
      RECT 7.130000 0.825000 7.300000 1.075000 ;
      RECT 7.130000 1.075000 7.800000 1.245000 ;
      RECT 7.130000 1.245000 7.300000 1.470000 ;
    LAYER mcon ;
      RECT 1.985000 0.765000 2.155000 0.935000 ;
      RECT 5.685000 0.765000 5.855000 0.935000 ;
    LAYER met1 ;
      RECT 1.925000 0.735000 2.215000 0.780000 ;
      RECT 1.925000 0.780000 5.915000 0.920000 ;
      RECT 1.925000 0.920000 2.215000 0.965000 ;
      RECT 5.625000 0.735000 5.915000 0.780000 ;
      RECT 5.625000 0.920000 5.915000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_2
END LIBRARY
