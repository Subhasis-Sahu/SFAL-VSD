# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nor4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.075000 1.805000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.075000 3.750000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.075000 5.685000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.810000 1.075000 8.655000 1.285000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 7.245000 0.905000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 2.195000 0.255000 2.525000 0.725000 ;
        RECT 3.035000 0.255000 3.365000 0.725000 ;
        RECT 4.395000 0.255000 4.725000 0.725000 ;
        RECT 5.235000 0.255000 5.565000 0.725000 ;
        RECT 6.075000 0.255000 6.405000 0.725000 ;
        RECT 6.115000 0.905000 6.465000 1.455000 ;
        RECT 6.115000 1.455000 7.205000 1.625000 ;
        RECT 6.115000 1.625000 6.365000 2.125000 ;
        RECT 6.915000 0.255000 7.245000 0.725000 ;
        RECT 6.955000 1.625000 7.205000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.740000 0.085000 ;
        RECT 0.175000  0.085000 0.345000 0.895000 ;
        RECT 1.015000  0.085000 1.185000 0.555000 ;
        RECT 1.855000  0.085000 2.025000 0.555000 ;
        RECT 2.695000  0.085000 2.865000 0.555000 ;
        RECT 3.535000  0.085000 4.225000 0.555000 ;
        RECT 4.895000  0.085000 5.065000 0.555000 ;
        RECT 5.735000  0.085000 5.905000 0.555000 ;
        RECT 6.575000  0.085000 6.745000 0.555000 ;
        RECT 7.415000  0.085000 7.585000 0.555000 ;
        RECT 8.355000  0.085000 8.585000 0.905000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.740000 2.805000 ;
        RECT 0.595000 1.795000 0.805000 2.635000 ;
        RECT 1.395000 1.795000 1.645000 2.635000 ;
        RECT 8.355000 1.455000 8.585000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 1.455000 2.065000 1.625000 ;
      RECT 0.095000 1.625000 0.425000 2.465000 ;
      RECT 0.975000 1.625000 1.225000 2.465000 ;
      RECT 1.815000 1.625000 2.065000 2.295000 ;
      RECT 1.815000 2.295000 3.745000 2.465000 ;
      RECT 2.235000 1.455000 5.525000 1.625000 ;
      RECT 2.235000 1.625000 2.485000 2.125000 ;
      RECT 2.655000 1.795000 2.905000 2.295000 ;
      RECT 3.075000 1.625000 3.325000 2.125000 ;
      RECT 3.495000 1.795000 3.745000 2.295000 ;
      RECT 4.015000 1.795000 4.265000 2.295000 ;
      RECT 4.015000 2.295000 7.625000 2.465000 ;
      RECT 4.435000 1.625000 4.685000 2.125000 ;
      RECT 4.855000 1.795000 5.105000 2.295000 ;
      RECT 5.275000 1.625000 5.525000 2.125000 ;
      RECT 5.695000 1.455000 5.945000 2.295000 ;
      RECT 6.535000 1.795000 6.785000 2.295000 ;
      RECT 6.635000 1.075000 7.640000 1.285000 ;
      RECT 7.375000 1.795000 7.625000 2.295000 ;
      RECT 7.470000 0.735000 8.185000 0.905000 ;
      RECT 7.470000 0.905000 7.640000 1.075000 ;
      RECT 7.470000 1.285000 7.640000 1.455000 ;
      RECT 7.470000 1.455000 8.185000 1.625000 ;
      RECT 7.810000 0.255000 8.185000 0.735000 ;
      RECT 7.850000 1.625000 8.185000 2.465000 ;
  END
END sky130_fd_sc_hd__nor4b_4
END LIBRARY
