# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.795000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.285000 0.305000  9.615000 0.735000 ;
        RECT  9.285000 0.735000 10.955000 0.905000 ;
        RECT  9.285000 1.505000 10.955000 1.675000 ;
        RECT  9.285000 1.675000  9.615000 2.395000 ;
        RECT 10.135000 0.305000 10.465000 0.735000 ;
        RECT 10.135000 1.675000 10.465000 2.395000 ;
        RECT 10.655000 0.905000 10.955000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535000 1.035000 4.025000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.255000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.085000 0.785000 3.255000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  1.975000  0.085000  2.305000 0.445000 ;
        RECT  3.765000  0.085000  3.965000 0.525000 ;
        RECT  5.725000  0.085000  6.095000 0.585000 ;
        RECT  7.750000  0.085000  8.120000 0.615000 ;
        RECT  8.925000  0.085000  9.095000 0.695000 ;
        RECT  9.795000  0.085000  9.965000 0.565000 ;
        RECT 10.635000  0.085000 10.805000 0.565000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.040000 2.805000 ;
        RECT  0.520000 2.135000  0.850000 2.635000 ;
        RECT  1.880000 2.245000  2.210000 2.635000 ;
        RECT  3.760000 2.165000  3.930000 2.635000 ;
        RECT  5.935000 1.835000  6.105000 2.635000 ;
        RECT  7.815000 2.135000  8.120000 2.635000 ;
        RECT  8.925000 1.625000  9.105000 2.635000 ;
        RECT  9.795000 1.845000  9.965000 2.635000 ;
        RECT 10.635000 1.845000 10.805000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000  0.345000 0.635000 ;
      RECT 0.175000 0.635000  0.810000 0.805000 ;
      RECT 0.180000 1.795000  0.845000 1.965000 ;
      RECT 0.180000 1.965000  0.350000 2.465000 ;
      RECT 0.615000 0.805000  0.810000 0.970000 ;
      RECT 0.615000 0.970000  0.845000 1.795000 ;
      RECT 1.015000 0.345000  1.245000 0.715000 ;
      RECT 1.020000 0.715000  1.245000 2.465000 ;
      RECT 1.435000 0.275000  1.805000 0.445000 ;
      RECT 1.435000 0.445000  1.605000 1.860000 ;
      RECT 1.435000 1.860000  3.250000 2.075000 ;
      RECT 1.435000 2.075000  1.710000 2.445000 ;
      RECT 2.120000 0.955000  2.465000 1.125000 ;
      RECT 2.120000 1.125000  2.290000 1.860000 ;
      RECT 2.695000 2.245000  3.590000 2.415000 ;
      RECT 2.820000 0.275000  3.595000 0.445000 ;
      RECT 3.080000 1.355000  3.275000 1.685000 ;
      RECT 3.080000 1.685000  3.250000 1.860000 ;
      RECT 3.420000 1.825000  4.385000 1.995000 ;
      RECT 3.420000 1.995000  3.590000 2.245000 ;
      RECT 3.425000 0.445000  3.595000 0.695000 ;
      RECT 3.425000 0.695000  4.385000 0.865000 ;
      RECT 4.215000 0.365000  4.565000 0.535000 ;
      RECT 4.215000 0.535000  4.385000 0.695000 ;
      RECT 4.215000 0.865000  4.385000 1.825000 ;
      RECT 4.215000 1.995000  4.385000 2.065000 ;
      RECT 4.215000 2.065000  4.450000 2.440000 ;
      RECT 4.555000 0.705000  5.135000 1.035000 ;
      RECT 4.555000 1.035000  4.795000 1.905000 ;
      RECT 4.695000 2.190000  5.765000 2.360000 ;
      RECT 4.735000 0.365000  5.475000 0.535000 ;
      RECT 4.985000 1.655000  5.425000 2.010000 ;
      RECT 5.305000 0.535000  5.475000 1.315000 ;
      RECT 5.305000 1.315000  6.105000 1.485000 ;
      RECT 5.595000 1.485000  6.105000 1.575000 ;
      RECT 5.595000 1.575000  5.765000 2.190000 ;
      RECT 5.645000 0.765000  6.445000 1.065000 ;
      RECT 5.645000 1.065000  5.815000 1.095000 ;
      RECT 5.935000 1.245000  6.105000 1.315000 ;
      RECT 6.275000 0.365000  6.735000 0.535000 ;
      RECT 6.275000 0.535000  6.445000 0.765000 ;
      RECT 6.275000 1.065000  6.445000 2.135000 ;
      RECT 6.275000 2.135000  6.525000 2.465000 ;
      RECT 6.615000 0.705000  7.165000 1.035000 ;
      RECT 6.615000 1.245000  6.805000 1.965000 ;
      RECT 6.750000 2.165000  7.635000 2.335000 ;
      RECT 6.965000 0.365000  7.505000 0.535000 ;
      RECT 6.975000 1.035000  7.165000 1.575000 ;
      RECT 6.975000 1.575000  7.295000 1.905000 ;
      RECT 7.335000 0.535000  7.505000 0.995000 ;
      RECT 7.335000 0.995000  8.400000 1.325000 ;
      RECT 7.335000 1.325000  7.635000 1.405000 ;
      RECT 7.465000 1.405000  7.635000 2.165000 ;
      RECT 7.805000 1.575000  8.755000 1.905000 ;
      RECT 8.390000 0.300000  8.750000 0.825000 ;
      RECT 8.470000 1.905000  8.755000 2.455000 ;
      RECT 8.570000 0.825000  8.750000 1.075000 ;
      RECT 8.570000 1.075000 10.485000 1.325000 ;
      RECT 8.570000 1.325000  8.755000 1.575000 ;
    LAYER mcon ;
      RECT 0.615000 1.785000 0.785000 1.955000 ;
      RECT 1.055000 0.765000 1.225000 0.935000 ;
      RECT 4.755000 0.765000 4.925000 0.935000 ;
      RECT 5.215000 1.785000 5.385000 1.955000 ;
      RECT 6.625000 0.765000 6.795000 0.935000 ;
      RECT 6.625000 1.785000 6.795000 1.955000 ;
    LAYER met1 ;
      RECT 0.555000 1.755000 0.845000 1.800000 ;
      RECT 0.555000 1.800000 6.855000 1.940000 ;
      RECT 0.555000 1.940000 0.845000 1.985000 ;
      RECT 0.995000 0.735000 1.285000 0.780000 ;
      RECT 0.995000 0.780000 6.855000 0.920000 ;
      RECT 0.995000 0.920000 1.285000 0.965000 ;
      RECT 4.695000 0.735000 4.985000 0.780000 ;
      RECT 4.695000 0.920000 4.985000 0.965000 ;
      RECT 5.155000 1.755000 5.445000 1.800000 ;
      RECT 5.155000 1.940000 5.445000 1.985000 ;
      RECT 6.565000 0.735000 6.855000 0.780000 ;
      RECT 6.565000 0.920000 6.855000 0.965000 ;
      RECT 6.565000 1.755000 6.855000 1.800000 ;
      RECT 6.565000 1.940000 6.855000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfxtp_4
END LIBRARY
