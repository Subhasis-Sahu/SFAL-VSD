# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__sdlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.850000 0.955000 1.190000 1.325000 ;
        RECT 0.880000 1.325000 1.190000 1.445000 ;
        RECT 0.880000 1.445000 1.235000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.530000 0.255000 6.815000 0.825000 ;
        RECT 6.530000 1.495000 6.815000 2.465000 ;
        RECT 6.645000 0.825000 6.815000 1.495000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.340000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.710000 0.955000 6.010000 1.265000 ;
        RECT 4.710000 1.265000 4.930000 1.325000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.515000  0.085000 0.845000 0.445000 ;
        RECT 2.665000  0.085000 3.010000 0.825000 ;
        RECT 4.080000  0.085000 4.410000 0.445000 ;
        RECT 5.505000  0.085000 6.360000 0.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.085000 1.835000 0.345000 2.635000 ;
        RECT 2.370000 2.075000 3.010000 2.635000 ;
        RECT 3.580000 2.255000 5.490000 2.635000 ;
        RECT 6.030000 2.255000 6.360000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.345000 0.615000 ;
      RECT 0.085000 0.615000 1.190000 0.785000 ;
      RECT 0.510000 0.785000 0.680000 1.460000 ;
      RECT 0.510000 1.460000 0.710000 1.755000 ;
      RECT 0.540000 1.755000 0.710000 2.125000 ;
      RECT 0.540000 2.125000 1.255000 2.465000 ;
      RECT 1.015000 0.255000 1.190000 0.615000 ;
      RECT 1.360000 0.255000 2.495000 0.535000 ;
      RECT 1.360000 0.705000 1.700000 1.205000 ;
      RECT 1.360000 1.205000 1.860000 1.325000 ;
      RECT 1.405000 1.325000 1.860000 1.955000 ;
      RECT 1.425000 2.125000 2.200000 2.465000 ;
      RECT 1.870000 0.705000 2.155000 1.035000 ;
      RECT 2.030000 1.205000 3.010000 1.375000 ;
      RECT 2.030000 1.375000 2.200000 2.125000 ;
      RECT 2.325000 0.535000 2.495000 0.995000 ;
      RECT 2.325000 0.995000 3.010000 1.205000 ;
      RECT 2.370000 1.575000 2.540000 1.635000 ;
      RECT 2.370000 1.635000 3.400000 1.905000 ;
      RECT 3.180000 0.255000 3.400000 1.635000 ;
      RECT 3.180000 1.905000 3.400000 1.915000 ;
      RECT 3.180000 1.915000 5.450000 2.085000 ;
      RECT 3.180000 2.085000 3.400000 2.465000 ;
      RECT 3.580000 0.255000 3.910000 0.765000 ;
      RECT 3.580000 0.765000 4.005000 0.935000 ;
      RECT 3.580000 0.935000 3.750000 1.575000 ;
      RECT 3.580000 1.575000 3.990000 1.745000 ;
      RECT 3.920000 1.105000 4.465000 1.275000 ;
      RECT 4.160000 1.275000 4.465000 1.495000 ;
      RECT 4.160000 1.495000 4.960000 1.745000 ;
      RECT 4.175000 0.615000 4.830000 0.785000 ;
      RECT 4.175000 0.785000 4.465000 1.105000 ;
      RECT 4.580000 0.255000 4.830000 0.615000 ;
      RECT 5.010000 0.255000 5.270000 0.615000 ;
      RECT 5.010000 0.615000 6.360000 0.785000 ;
      RECT 5.140000 1.435000 5.610000 1.605000 ;
      RECT 5.140000 1.605000 5.450000 1.915000 ;
      RECT 5.660000 1.775000 6.360000 2.085000 ;
      RECT 5.660000 2.085000 5.830000 2.465000 ;
      RECT 5.780000 1.435000 6.360000 1.775000 ;
      RECT 6.190000 0.785000 6.360000 0.995000 ;
      RECT 6.190000 0.995000 6.460000 1.325000 ;
      RECT 6.190000 1.325000 6.360000 1.435000 ;
    LAYER mcon ;
      RECT 1.525000 1.445000 1.695000 1.615000 ;
      RECT 1.985000 0.765000 2.155000 0.935000 ;
      RECT 3.835000 0.765000 4.005000 0.935000 ;
      RECT 4.295000 1.445000 4.465000 1.615000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.525000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 1.925000 0.735000 2.215000 0.780000 ;
      RECT 1.925000 0.780000 4.065000 0.920000 ;
      RECT 1.925000 0.920000 2.215000 0.965000 ;
      RECT 3.775000 0.735000 4.065000 0.780000 ;
      RECT 3.775000 0.920000 4.065000 0.965000 ;
      RECT 4.235000 1.415000 4.525000 1.460000 ;
      RECT 4.235000 1.600000 4.525000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_1
END LIBRARY
