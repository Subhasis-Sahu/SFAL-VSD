# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__xnor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.255000 1.075000 2.705000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 0.960000 1.285000 ;
        RECT 0.790000 1.285000 0.960000 1.445000 ;
        RECT 0.790000 1.445000 3.100000 1.615000 ;
        RECT 2.930000 1.075000 3.955000 1.285000 ;
        RECT 2.930000 1.285000 3.100000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.913000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.795000 5.295000 1.965000 ;
        RECT 3.725000 1.965000 3.935000 2.125000 ;
        RECT 4.585000 0.305000 5.895000 0.475000 ;
        RECT 5.045000 1.415000 5.895000 1.625000 ;
        RECT 5.045000 1.625000 5.295000 1.795000 ;
        RECT 5.045000 1.965000 5.295000 2.125000 ;
        RECT 5.505000 0.475000 5.895000 1.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 1.450000  0.085000 1.620000 0.555000 ;
        RECT 2.430000  0.085000 2.600000 0.905000 ;
        RECT 3.270000  0.085000 3.440000 0.555000 ;
        RECT 4.145000  0.085000 4.315000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.570000 2.135000 0.820000 2.635000 ;
        RECT 1.410000 2.135000 1.660000 2.635000 ;
        RECT 2.810000 2.135000 3.060000 2.635000 ;
        RECT 4.625000 2.135000 4.875000 2.635000 ;
        RECT 5.465000 1.795000 5.895000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.645000 0.860000 0.895000 ;
      RECT 0.085000 0.895000 0.315000 1.785000 ;
      RECT 0.085000 1.785000 3.480000 1.955000 ;
      RECT 0.085000 1.955000 2.080000 1.965000 ;
      RECT 0.085000 1.965000 0.400000 2.465000 ;
      RECT 0.105000 0.255000 1.280000 0.475000 ;
      RECT 0.990000 1.965000 1.240000 2.465000 ;
      RECT 1.030000 0.475000 1.280000 0.725000 ;
      RECT 1.030000 0.725000 2.120000 0.905000 ;
      RECT 1.790000 0.255000 2.120000 0.725000 ;
      RECT 1.830000 1.965000 2.080000 2.465000 ;
      RECT 2.390000 2.125000 2.640000 2.465000 ;
      RECT 2.770000 0.255000 3.100000 0.725000 ;
      RECT 2.770000 0.725000 5.335000 0.905000 ;
      RECT 3.230000 2.125000 3.555000 2.295000 ;
      RECT 3.230000 2.295000 4.355000 2.465000 ;
      RECT 3.310000 1.455000 4.805000 1.625000 ;
      RECT 3.310000 1.625000 3.480000 1.785000 ;
      RECT 3.610000 0.255000 3.975000 0.725000 ;
      RECT 4.105000 2.135000 4.355000 2.295000 ;
      RECT 4.635000 1.075000 5.295000 1.245000 ;
      RECT 4.635000 1.245000 4.805000 1.455000 ;
      RECT 5.005000 0.645000 5.335000 0.725000 ;
    LAYER mcon ;
      RECT 2.465000 2.125000 2.635000 2.295000 ;
      RECT 3.385000 2.125000 3.555000 2.295000 ;
    LAYER met1 ;
      RECT 2.405000 2.095000 2.695000 2.140000 ;
      RECT 2.405000 2.140000 3.615000 2.280000 ;
      RECT 2.405000 2.280000 2.695000 2.325000 ;
      RECT 3.325000 2.095000 3.615000 2.140000 ;
      RECT 3.325000 2.280000 3.615000 2.325000 ;
  END
END sky130_fd_sc_hd__xnor2_2
END LIBRARY
