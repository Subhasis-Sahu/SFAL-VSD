# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a2bb2o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.075000 3.645000 1.325000 ;
        RECT 3.475000 1.325000 3.645000 1.445000 ;
        RECT 3.475000 1.445000 4.965000 1.615000 ;
        RECT 4.605000 1.075000 4.965000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 4.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.445000 ;
        RECT 0.085000 1.445000 1.685000 1.615000 ;
        RECT 1.515000 1.075000 1.895000 1.245000 ;
        RECT 1.515000 1.245000 1.685000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.075000 1.345000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.275000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.920000 0.905000 ;
        RECT 5.275000 1.785000 6.365000 1.955000 ;
        RECT 5.275000 1.955000 5.525000 2.465000 ;
        RECT 6.075000 0.275000 6.405000 0.725000 ;
        RECT 6.115000 1.415000 6.920000 1.655000 ;
        RECT 6.115000 1.655000 6.365000 1.785000 ;
        RECT 6.115000 1.955000 6.365000 2.465000 ;
        RECT 6.610000 0.905000 6.920000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.360000 0.085000 ;
        RECT 0.175000  0.085000 0.345000 0.895000 ;
        RECT 1.855000  0.085000 2.025000 0.555000 ;
        RECT 2.695000  0.085000 3.385000 0.555000 ;
        RECT 4.055000  0.085000 4.225000 0.555000 ;
        RECT 4.895000  0.085000 5.065000 0.895000 ;
        RECT 5.735000  0.085000 5.905000 0.555000 ;
        RECT 6.575000  0.085000 6.745000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.555000 2.125000 0.805000 2.635000 ;
        RECT 1.395000 2.125000 1.645000 2.635000 ;
        RECT 3.175000 2.135000 3.425000 2.635000 ;
        RECT 4.855000 1.795000 5.105000 2.635000 ;
        RECT 5.695000 2.165000 5.945000 2.635000 ;
        RECT 6.535000 1.825000 6.785000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.135000 1.785000 2.065000 1.955000 ;
      RECT 0.135000 1.955000 0.385000 2.465000 ;
      RECT 0.515000 0.255000 1.685000 0.475000 ;
      RECT 0.515000 0.475000 0.765000 0.905000 ;
      RECT 0.935000 0.645000 1.270000 0.735000 ;
      RECT 0.935000 0.735000 2.525000 0.905000 ;
      RECT 0.975000 1.955000 1.225000 2.465000 ;
      RECT 1.815000 1.955000 2.065000 2.295000 ;
      RECT 1.815000 2.295000 2.905000 2.465000 ;
      RECT 1.855000 1.455000 2.065000 1.785000 ;
      RECT 2.195000 0.255000 2.525000 0.735000 ;
      RECT 2.235000 0.905000 2.445000 1.415000 ;
      RECT 2.235000 1.415000 2.620000 1.965000 ;
      RECT 2.235000 1.965000 2.485000 2.125000 ;
      RECT 2.615000 1.075000 3.145000 1.245000 ;
      RECT 2.655000 2.135000 2.905000 2.295000 ;
      RECT 2.955000 0.725000 4.725000 0.905000 ;
      RECT 2.955000 0.905000 3.145000 1.075000 ;
      RECT 2.955000 1.245000 3.145000 1.495000 ;
      RECT 2.955000 1.495000 3.305000 1.665000 ;
      RECT 3.135000 1.665000 3.305000 1.785000 ;
      RECT 3.135000 1.785000 4.265000 1.965000 ;
      RECT 3.555000 0.255000 3.885000 0.725000 ;
      RECT 3.595000 2.135000 3.845000 2.295000 ;
      RECT 3.595000 2.295000 4.685000 2.465000 ;
      RECT 4.015000 1.965000 4.265000 2.125000 ;
      RECT 4.395000 0.255000 4.725000 0.725000 ;
      RECT 4.435000 1.785000 4.685000 2.295000 ;
      RECT 5.135000 1.075000 6.440000 1.245000 ;
      RECT 5.135000 1.245000 5.460000 1.615000 ;
    LAYER mcon ;
      RECT 2.450000 1.445000 2.620000 1.615000 ;
      RECT 5.230000 1.445000 5.400000 1.615000 ;
    LAYER met1 ;
      RECT 2.390000 1.415000 2.680000 1.460000 ;
      RECT 2.390000 1.460000 5.460000 1.600000 ;
      RECT 2.390000 1.600000 2.680000 1.645000 ;
      RECT 5.170000 1.415000 5.460000 1.460000 ;
      RECT 5.170000 1.600000 5.460000 1.645000 ;
  END
END sky130_fd_sc_hd__a2bb2o_4
END LIBRARY
